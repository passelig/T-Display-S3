PK   U�tWm扴u  �    cirkitFile.json�]Y�7��+:歋�����L��R��I��e1�E��l�^�~����M�f�Jv�lŮ��j@"������m�_�jQ�7n��l����ʻ��|S}�Ͽ%w���j�[/~��g������G���O��[�,/dQ1��B�L����Rɕ5���1� ��wC��+�5ɘ�e&D�<g,#��NXS��.��nhlU;�
K3%�̄%<�55�&'Ԗ��ap0�k�� �&�Y�kbK��3��	���jg2UJ�8/9�
�^3sd�8S2/��*)���~�֙Q&�W��n���1\F�vF�\��Һ΄+�̔y�QW�\��p�D��%/�����Lm��q�1���/�4��m��p9� �Q[�q[ep�-n8%��1qT�R&�_w�GRd�u�\���$�\�f�LM�QSǄ
hj��Z`����cR4�BM��uljUZQ�23��r�,M��<�b\rWiF%��Nq�n8��ë4T3��
а�h�\ᙁf����3�6�^@��f@+�fF=sl�K[�J��Y��j�啧����4-4QrD����ehx\�mqĲ��=��@��q�>ꙇ�
�2�k�M����Q6!�	Q���>r�`�4Fm��hJc����)��:&��4f� 4�1S�tД�LU^���.�|a�'�Ҹ��������l�D�W���8l|<�o�Ч�)�bu&�7q+�GV#�RQ������D��1]4g��8��b�T��$kg3]�گ��tQW
�6��ԑ�)'��F�1@��h�#�=��Q�j�P>�D
�t!M�/�{�r��� ��f������н��[B��A�*ڱ�b*<P��.,���?Q���"��.��*jO�*�BP�I��$�b�P�$�=z)!�]�|���p2|��ʉ�_U����� ����X��**f����H@�%�§�@�
��/4�?�
�!�q^���q^���q�	��qh�;:�D�P�8��T&�4>=�����q7�����D�ǒ+�!Yϋ#�Dt4�:��� k*lJYCæ�W��`渦��%�54�8�����xI�4����
ILAf�?�S�Qi�L�(�`c
2v��W$�f�� �K�6fJŁCf)4�䑂�Ʒ�_hlj�h�����v��6d�rO�M��ᩰ$Tx*"	���JBE'�b�P�iP��i�K�����/M`��t�А���vCCFx*���L�8d��2�8d��2�8d��2�8d������s�L�2�SI����CFx*�x����T&�.8d��2�b�!#<�I#2J��D�K��i�2J@&���;x�(�4裓>
<d�@^�A1K$=�lx�fi��xL�����6�CFx*�|������-��o�{q7��ܸ���!/]�X��M�6��w�M����7����0eV(j3)��;�������d5�|��[�\�O�I�j2�_>���0S�rQjjTnEM�Bxf�28�u�ޥ�<�L��y�{�y?�PF���ɯ�4��ѧM��Y�p�����M�)���%H��45åy���d�����N��Mu�l-Df#�p��L�{�F%��i�X�_Cc��W*���U�
hj�fG���:45J�F��vU!�(3��b�ʺ�5ϤVRp�tY��g�� ^>3�l�L�X�!�rŝ�*�[�U��)���-��w(���3�2� 3GW�pƼ�$YA���e-�\	�Յ!���(�YfчM�R�у�e(D�	hjԙ�
Q���<x��(�U���s8y��҇��I��\��k�%/�������
��33�}���BTEĹ�\+�5)JKc:�4����d3u�\����;b��Kob��]CS�C�a �s�a/��aoԯaS�a�c$
�HRr�/��.�5���0����E���������W��i������n|�|�;�avثG<�H<ػ<��&��d�A��A�)
�c9�� x�Rp9	�S����4 ��D$"��� ����������?�������&)��$s �6� ��Uu�M�	�`�
�`�p��1�s�N5��b B��x��h  E��$�8���T))8�jF<�z���Ab"�9� ����$A�Y��B�9��D�9�fF�9�j�&yR��"]
� 2��4!��xm���H�ǔ�m�!��(Bs��h�*	�^/㍴ȅL�%` �@Q~� �k� XOX�7�-�s��`�s��.�s�M��s��+�s�M���Y�x�i��"'�j"45u��[d��@&�� ���g ��:.�n���_dk� ��7�n3��et��Z<��Z<�)�X\�_��m�� m��9@ۦhж)��m�� &��-�� w�&��x��(�$��U�d��9�j��&9�W3P���x��	`�L��s����ֺA���z�l~��,�TO�թ������GFBY��e�-JO��P
�O��X�\,�	�;���ܺ����-�&J��a��4��r�E�oj���e���L�fK��}zȼ�=ԟf 8�o��Z�3�!���xp)��jFd5��}�\D����øW��q.w�!����rM .���� w���ď�\3~�܁�W#fE�+�w�a�p����;�0���3�A	Z'3~@�G,p����� ���!�;p��9��hs������>
Yhhb�IG��~>�������"��F� x�|����*l����3`����#�K� `���~>�;p!����͞�,�����!��g��f��z	P�<U|���8��Z4Xs*(7ԼE�TJ�A����~ ďz�@\�� ��� q Z &v��� �!�~�1ٛr!X ���}i #���&���P�[���z��l� 䴜�G�i2Vn��7��o�k�xypl@e��Dc$�&!\#��#$�l`�
�E �!ăDB;��DpMɾ6~�$�a�~�ń���- � [-��3s���}���b�}Gp���؏M �A�c�^ܠ+4��Jn�E���07������ �EP��'�a�r�ɗ �+<[������=#�������	��ӤM��dM��dM�����BSc�w�豍�I����Ӱ~;4�~?4�~�84�~�<4�>�ǹh2z���g����/~��E�qyU��M(Y���.@П~��.���'��<+J)���ՄJ�������������ջ���g����.x�4_�ݬ�f�t�;��q�8��nw����$��S�Z�f��O��_���C�O���d��~\~��wOwv_�[��n��r�,�黍�ϧ��yr���Ƨ|�T���i�d�8�v���\�]N<+���r�\�ux��Ka�5�.cD΅T�H���������\�+/դn"֛����o�iι���X���|U�ǀb&w��f�w+��2{z�_��M����NX=��Q-�m��;�	5��%b�k�&��k��&���s�}� ��g"t����HE�\+���7�M��	�}��D��P�0C"�����8Qv��<<�$s�9�`D��,=qr�ǔ��ϬxX$è���V*�T�R:P�p�����X:(aϧ��i�]�Y8�@��ٓ�\�v�5��X����h �����S�\��6�=��fΙSX���~���w�+�?=���i�^LP6��_��b��c�\NМ�^e��Y������+��L��z	���	H� '���0���������-TϛSt8�l���#�=��0�!�M1y$��滌r�U蛫!�5�ƫ��0��/��s&5g�c��q%��]�3#M��2��Y�mn�)+�嶧@a�.����UYL��,�|��sC��Ak� -=j<��O����u �[�D�� �x ddn�:�A/kj�#��+�*���T�CG/��7.��Q\�)V�`�f�\xL�Ċ�ֈLi������i�EP5V�9��[K�+f�{�[�	�T��t/GZ%({)bD(��M�����눹=���!޲=ijI[��A�Z%�/CFZ67�//?)/X��x����s�\Ƌ�e��*�s^(��M�dö������x�6X��F>~�����!�
��oU^o���o�_UOa����7s�	U��4P��q��� �&��ҟά�>HV�q�-L�y'_Tq%i�-t��@rDȠbh�����d�gs�(/�G{Q4�s�C�DH�x����R8S��Y.Y�	呯E��,�u)J�W�
(1rP�^�ۖ�!d@t��EF�Ly���z�TyCP3�VZ��w��B�6eD������3]y7��Z+z����]�&���asyս���߬V��X�����<4\���S�m�=�
���%�s<7��f�81�6��Դ_����b����qj�/ȱi`INM�E96<䩩�0'��ǡw��M�u>�R��h
k�"]���.��?S��)H���8�tR������� ��ڠ��~�W��t(rg	�ԋv�=T���p7�����t��D��^�L�%��p"�M��7P�WdN��5���Y���H��B�[O�����p�o���|����(ݾg\��w�N���J�F���iK{�RK)UV�9ψp:�2����B�����u�t�[W�m��|�K���v��<x��4�	��7 �`,hA�@����m�>�t��6u�t\Ե_�YF�w5������3Մ��"~^V���;k�\޼���5l��һ�R2.����C>�\��GW}w��}�q���?/���i0�����<�7�g��g���y�~v��{�f�v���j�^�~�s�j�,�!��?���5O�o�{\/W����cC���������mh������w�gs�zu��mk�q~�����ع�}���C�>|y?��!�u��b�Z฀�뀃[��n�4e/�v
��v�C_F�C���:%�H:9DC�$�C4	�Z!��/��|�'�r�t���u����k����QR�nBv��!X�����:��H�a��uA�N	5	�����P�P�]�݅P{N�:`���u�N+:��u��,�ࠔ��_�����~_�`o��.��B�ٕs���t�[U�TJp�t�(58TRQ�������� ��UD��v��{��n뽳��H��m�w�^mp�U�MOVMu�%ua��.A����	���qw�ವO�����^bP����;�����5��,��pK�,p�.��6m�p�Иv@�2��zT'�fa�ʋPv��O���6e��v
epw!ʦ�)����Lۺ�vc]A�F^�p\��낣c���x���k��
8�cU�Ը��V[!�q��ጛS6]�"�c�@{�@����Av�"$��P"D��an
��`�5R߷���ػ�	;����O���%!���z�
j垁���fd��QR�����)���<^��������1�u{�i��;`7(���]�4�DE:���HI�&_�����Q�uz� iҾ�iu���I��3���F8�p{�"�U� ��N�[ ����E�3�.)�X:�]���TH{Q<��N�(�:�n�4	�Ӻ����?I��a�0pq�oz	o���"���d��:�n�4�ӺݠH��?T����%�Q�xK��] v����n����I�n�q�̡���_Bx\��po���l�A��v�Ɔª#�Ά^���n��d�b�ݤ�ᔳ޾��Q�ίC��m��e��m��!/Lگ˝��{��[ү�ڦ���Kػ<�Ԇv�$u���nލ[><������f�?lg�X����\��|��?|�����}چg��e��PK   �rmW�\>& %& /   images/27abb4c4-9cc3-40d1-807d-7d8b935f4094.png >@���PNG

   IHDR   �     @o�   sRGB ���   gAMA  ���a   	pHYs  �  ��o�d  ��IDATx^���_�u����}%�z�B	�@��b\ �v�S�'�ɓ��4'N\�c;�-6cL3��E�{o���>��ܻZ�j�����럳;�;wʙ3gΜ93w�܂={��������G�0������h���������((p0�@��{Ba�w�+(:����o῅ �������رs[�tF�(*,,��D��
�:���4��D2�#���~�c�QT\�I��STX�
+**��Ύ(ֵ��P銢��[y�H_��(..Q�Pxw���5^R�=]��Gt�с�H�t�"ߋV���}Ƣ������.�����,O�h�
k\y�$i����Wf��]�� �M	uI~ht&nM�n�DwY����~P89�JJ+�Pt�w�*�0���/��c��jT���"� �O:1��)�%�jX��H�Mm�0<�rlA�J2B+�'�z��T���"�@����-���I(|Y��R ��]�U�����Q>	 �;��Z��`S/%NuA���"yJW���XT��$��T���%��\� ��BաH�������L��Ӷ�wcX�bu��Du B�NW(Ĕ�H�鎪{����GIaO�w�+A��1���w�U5\�8��o����m7���jy	�ڥ�C�g���9=���~it����Z��0�GP���A�o�`5y���F���W���_��P�ki�4�ʴ�V��Xx�1u�Ə�C���@ք%tC��OZ�0>��M^��~��d���9�S,�)�����Tg�t*-#�+}'��}��X�2[ڻ�U�h���c�رqU45�W��Y� �=t(`�N]�7�PYQ��艮���PT���"N�69�ϟc'L���*�}��
��u���X�u3��EqY��*	��[*� ��d>X �h����&si���i8y$i#�3nکq�Yg	��A�ς!�A//C,B�ko�G�ʴ0s���!<�A�ih�8+�� )i��U�ƴHø�}!����@S�2��A�3���4u���~�طg���'�k��nА��u*��Dϲe�c�����y"	8A�ND}�#�\*�c�h�0����Ғ�(�(W)�Q���ß�d���"'N� oް6����a�W��ikj������(��%��]�b��C��-&�h�D(:%�4d�����v�wD�4R����9sc���jxM�&�2L�����I:R(�ie�-�x� �+��Oc��"�ЖXH'H"K�T�hF���
��V"锤5n3�jc��pGǒ�)oO�z��x�5QW7"J+�c�έ1fhEL�q�ҔپV_�g�{!�,z.::Z��#F��~ܩT���)	?��_����XfY]mu>2�uݻb��W׉�*�;�o�����mҲ;�o��;��������3�̲�ߣ�ʪrk�nۡj[ia�k`4U �3m1���q��)@�UB_�FD�yh�adV� �"\؏��T�����+��]X�@��N�>�� ��V��MY��%�*ѡXL��\)/�SL�-K�c��M��+�ƀ�âBc{Ye������7ƤICb���)��~�م���ϊOm��>2�@�AGOO�n���lax�z3aZ@㱣�'>��q�%'^��ί`Pþ��ꫯǺM;��]ڷ�S1)~�ӟ��|�;��(����M7�����ֶv�]6:e*�K붶�+/�jpԏ�SB�fa�^'ڲS��O1'ڻ:�)iL�k�h1ū��Q:�	��x�J�ӭ���m���h�f�5^�2)'�(�)�z�%tL�����t�lQGuA�TJv���n�Qc�FkK{l޸>v�����bĘ�u�vѬ�^C?ue"ٮzcR��N��!~u�O�ߡ{]ʔ������)Lu��-�-�}�i޽�1Z��	��?��?����k������]wF}33�B����g��nx�yԨQ1eʔ�7o���a�a��عs�����$ �3��7!Ǝ�wﰩ�D�����ڄ{Kk�y{i�77EUum��q��hm�U��H9�Nu�-�D��]�ˤ5YR���ݻ����K�+�g{��~�ھE4��m���~�i��d@`�k1�$D��v���c��u�X���Lei�?6n�!u���%���]ӯ����G�6^̯�k��&��N-�N����1�p�L�S^	1t$��S|�+�Ǐg�9�'N� �6����[��;c����W�Wq�i�Y#�u�'N�~�7b�޽�Cbr�$�1z�X��f�[���4k���#��>D�i�5�j"����GKK���	�c��x�ǥm:c���J�W�����K�ūK+oA2L�Q�����G~+V�u��ǀAc떍�ܓ�ǫ�-U��[7�5k����+���)�R'*5ݭ-M���%���c����v��ذn����z}{�4nW{�F��4hhT���IK�6z5r���[��Y�.6oZ���ŵ�
�L(��~x$p��1���z�̀��o�5��q�I1眹)��	5!���!����SN�@&{09����s�=��ܤ}qI�W�%t�+�wt���&����ε��_e76�D��n�Y��gO}46�hdװ�,zp��%1~�h�.�ilۼ^
M��,^$�\�����!#b�m��OĪ�cЈ�1k�Eq���bƙ󣭠_<������/k���ƫ//��/��2�c��gɆ� &Θ��������_f�aCGƖ��ٺ?F��qcj�I���M�cذ6��1���e���*����d�vI��3�AqJG���%��y������ĺBVw��	�$��a��s�ICR.�}!⚚�8��S��J� 6��Px�� ���2.�h_��^�W��Ǵ��h9����)�G �CH1!F��N9U�¾X�|Y���Ķm[��%/Ee�8}�̨�y�]���51i�)���y1cꘘ4~p�1kj�����)k��P�i�v^o��zTVT�<�P��2%�Nsgψ_����k��Ǝm�c�=~J4���K�.�^x!���#GO�!ÆK�ާ�f+P9���tB��z"Ȭ�������?Vd
�eD34�I2%�,A����N� 炄X]Um�� A<��Dyy�Cz�Fr�$�=�|�&\�]��ÐI2�µ{�˕\�5ߩ	�-Ě,2�f���H��S'O�!��ěo�/��t,|��h��1��sb�AQ�_lܴIګ$�O��j떖f�o������kd�;�b	Q�̄���aL�<5�mJ���,��%F��'����%��ԉ�b���8���c�isb�ɳc���Ÿ	�ă4!C�v�-3P����:lVc���mR ��Ǹ�gŐQ�I��)k��]�PWLg�"�wI�D`]h�n����_Ҽ��bnOZ�I�mGZ��ٵ�Q��k�D���\����Pv�1O���6�k'N80���+�ӳu���V��I'͐檊�}1�^�>N>��7n�ҵGCcc4�.U��Q^U�����U�e��o��(�����E�sc��-a��K}�J��?�3�P�읻�D���"��VC*ch��(�jsxf���y�Fu���d�=�()� ި~���]z�5q��>�����n������is������S^����n��G��`��D��o�>ٕ���Yw��9 ��e�1~�d_�$L:Rà�%�ʤy���K%�A7��4�\�l�̵J�y�Y�mKX:%<,�b������6��Gr��!1v�D�+�*��5�A˷Ȥh�]%�a#��6��+����.���^�<�X<��ӱk�.�NusY��M�����O���p���~t0��O������h"�̓:��N/�H���f�Qq�%�ǸQ�<	d��[�ݯ�'n�Ἐs�eQXR-a�y�%<����N0�P�)�b*�{[5\�y睱u�V�	��{�ڲys�uƬ�:e�N&���ͧ�t$� Ɠ�S��'J�%J�p"�nh5r��@��Z;�$�m�,��zn݀�(U�8��Y����UVZ!��*\�Hd=6�Ϝ�N;7ʫ	k�]Q^Q�a���D����v�'��%%*C&��G�!et�P'�32�#��D¼Ru�6��dm9�Z��9�j2\V�	k�l�11l��4hH�����[��ysN����9��E�ῇ�X֟'Vb
O�^|����׿{��P1��c��$8+W���o�;v���Ϗ�Ꚅ�\��L0��HjT�%)͒ve1�r/3Ca�))f';ƒ	�C����@+" ��h.���j0�׸j<^4�V�����>6�^��{��#������qc�(e@[C���X�rU�ݹ��yО;wn���6�?���e�hc
�����TO�h�d��#fbo�f�f쁘(�z�������5�#��e�UXe�#��w=�_!JKk����	`�"F'ӡ ��G�ٿ��X�h�����$�%�o��VlQc�EC}��`��5/�� k&ٽj�����K���W�,Ԍ~a���b?�����lg�����a劥������W�7�Ǝ-�P�_��4�SF:�ht��C9�;QZvp,{��x�Ņ�n�۞��]�f,Y�l�޵-
�؋\C��A��ƶm������W8�ވ���M�Ѝ;>�kk<R�D�M�ʔI6������~�)��$?D��2�-�aäi+ʢ���t]��L`q�L�Z[Z�F#�Au�%0���A�� N��$�{�O�^���a�\��۱f��رc{��g��ҥ˽�Y_�[�&���[�k�ǆ+��v�� ?�~��!Æ:ݎ�;c��ؼyG�ܱ7�m��w�Q����ojج�M;Ϋ��Ф�歱Ei�l��6oQӕĈ�#uM�|���-[�
G?i��:#��b����i��ظnC�Y�*V�^#����i�O�����������3�n�֯��k�J��hn��'N���8C�N���� 	��Jڛ���z =J�,����IV�(��ₘ8vT6L�Zg����\�KAꈝ-�aݦ�ׯ:V�\�6n��G����0g�>#f�:*N(���<[7o�O|��ؾ�QLC�a���N:9Οw^,_��l�vٻ��
��S�%��k�3f���8V�^��Ip�/��8i�8�䓽�W�ْ�	4������QSQo�Y�U�b䈡�,��s�~i3&��3o�U�~�jbP]��I�՚��c�:D���aC�;�{	��:��S��wˮ���연t��,��kc�:	O�R��JAs�F
�jb�.�R��4���N�����EL!4!Z���NC;���}AƵ+�P�$t^��_��'O�g�>;
˪V�WۯV�Bu�z�a��'?��L��Q\N�J�t�o}�#��?%'N� oC��ñm�^�4%����:tX���e�vǲזG����MC�]Q7hhԔw�ӏ?���k��0�FL�Sf��3N���5�&�ċ�	����V,mE)�g����#�07g�Lo��t2$H��V<
���]gģ�AQ"!F�1�Sy� ��a�Ȇ�u�'��M)���Nr�0K��6�	��;b���e:��Ҳ�$��4�2N;��<x�M�
u�r6��t�1cF�Ï<�}�ť�Q"b�H%Tq�����r"�
�����O��Ob��}jp��ɗ��$N?��8��Sc��ͱk�>](�b���I[l޴JC�1��k�T�P�� �?*&��7rqiZǤ�)�F�<���l�&	7E(-+
\š�	&oP�y��wބӯ�Y]@+�=��7��G�i�╏"�d�X���4�fᕐ�^�K+�yLH���� �
�H靺.�K{�����&�M?�]�Ý:�!��2	'u)���N�	c���7�Z�֭�R�������Ko�ܳb��	��D�	���x�%ָ�z�
`�b���]e��1���53l���u��hioQc��4�B���b5Ba�k��Z0�9;��s�&����Z>$�J�	�����+�D�xTBf!E���#��X�III �T��ˠ8��#�!�Y.Wqt
cNȌ��T_y������mR��>ȟ�A=�{xNEB_0�Xge�]yt8�R_aQ��6bdTUWω�"��MѰg{lX�zl۲6���bb��ZY��Bm f��`�(D�=����^�������42JPڮ���H�Ӑ!;����ȟT�ᔰ�)�����N$����c����s�ʑ�p�8�#$�˛4�����׏N�(d��T~�nr��D醺Au��xO��r՝> ���GC���j��tD��Zȯz+��!�邏��� 77Ի�y����k���bڬs����yN$��)���_�2V���w�GSKO�rc�Jd>X�H�Z���,LF�	�nn�fMv�bj��N�@���9G�3��OP�&&���'S*�3^�fl_0y�f: 48���H�O�DH��y�@im�C'x���'�3��f�˙
g��2��M�Q��ċ0�F�P�'��� ݕ�v��d��塬4r�V�b���ޮ<f��E�ڃ��p诼�4f͘��:=.����o�0�?�pBx��m�����X�zk�o��fL�dF$a���b�.jE�ʮ)����N��V��hR���S�!n|�?$Her�`��	16�y�>K�HH΁��=��0�!�H,&H��*֓J�9�M",�}2�(xB����<��0#�TR:Y�6�PYt_T��q�O^��l��V]�:�B���h%=���+/97���ߌ��#��D�	�=;7����ǒ�b�&g޴"Mh�350O!.���OB����Y��8���$�?��B��J�Oj��ο,��&o�Jn��r���]@OS>��:����o���xRF]�a���x'QxZ5����iOWL��H�(K�����N:=#adP��$e��%�iΏ�b"�)�6p@|�}W����`�4�iO$��_7��4Ek��`ט�Z`�Sa����R������[�s��.��NLw�!5Dj0����OCo��p�^Fx�	��q���&:f;�$�+�|�e'zL3y�OW����\�
��t9��=���=k��������u)-�Ht�$Q�.ʏ_׬��|��$�2S��e<q<\�&FX�_Cc���� 'D�[�4��1(��I�X�DVb�����֏�⸓#m6�fD�K")Ș�&IW�3�FVC�A���m��F��x�G�-�,�ՠ2X���(�s����3!��@F/	�X�W�����H��'��)�P�^�YZ�u ��9*���p�_�}s�4s��g��W��-�t�U'N� ��WEu�a�
_��� �	����&I�OBlF��)<5�b�1���5ȁ{a��p��r)]j�\`�߱YcC���Wʛ4��?|���	:R_�%���@�,	�WG2S�@�RS�r3�������'�)�3��O2�_�He�|J���)E�l�$��9}'N� �?-N=�L5
��ր���U1���a������z���H��y�<���$��>�')H�P^�AZ�q	WJ�:i=�Jpi*�W�SRj�#B��T�x7��ʤl�[�x��f��}�Ҹl�Vl�esڒ�Ax��M�Y�U��n�P��t����Nᩩ�uCG:�D�;!PS]c����&3@�0����`�L� �61;��h~�;�'iy5Hf�ڿ����X�P�,�xsA�!%�nR�ۑW�P&��EfI~��4PgӧH�Ul��X��!^�R|�,�_��S�l$>��tU:�RQΗ��D�0��b�i��R��U*��ښ��j�>��q�}�����`cvS#'�HB�+
�əMS�>'=���>�Y���9��������>K�\��~{���H� 
�X��|Y?F�R$�, �C	���)q��`���:�9��4�])�V�fQ8S*O��Q�y�S Q��L���CW��T���Go�.>��'a�-��	����2��ˣ�4G�+������������ *u<����g����{-�5&�60!JZX��q�g������f��g�ٛ�M���>�˒ٟ��*���N��e�euª?#Q*�u�]�;aFOV~��yB'Hefa�[Z���zs�J�y��kH��Fs��<
��hB]RP���BӮ���uv ��/}h��f����&	Pf�$��e����TVDOE�6���Ep,��xK�z��.�{8@�ڇ���>=��
����c�x�����n�>�^�z�mhJ,*0'X"gT1���8�8���a����A&�fH�KS���+���� �y�;�nx|�Ո��/�3@�AZ�RFJO)�AsAE�B��R�й;*8+*%&�3*OH� ?���!=�Q�ȃ�d��ȼ@(A�[}ī��(̫��O�B7�

e&H�'%	�xk$������YW-8+>��y8��?$bΙ�k�`���Y�,
�)l����e�����*���� H�������?���`�PՐ�~�73O?���L�0!����,���(v���W��E��O������Ly���ћ��g^x#�6��%�Nm�XlE� ��*��Pacs�
tE���)rCf��-/^���Oa@1��p�	�Q9<jBf��ߩ��2o���������6�'arB�(IƏ4�d�!�%I*��3��\%���~6�6�� �V���\٭��Q(�ڢn��h/:)v�xF�Y�X-�«%���+�����=�����=��hQ@�E��k�}�^��sX������7�qхQP*��
��bD߻������������������#�|D����@[@Og��}v�>��R���O��O>�F�����;�������s�%���=�yO�s�9q��׾�5����x��|��i��L�hD�>��V�4��ъ��44�V\T�<2%���g�8��a�eaa��e�,��f�!P�ƨ����ˢH����2��#�h�c��p8��5�)*.�5�8
�+�6t-�HRXD:��*Eo�d,��V&�%r��)�Tr���"�E�BQ�ù��
_TZ%e\��t�3��Q����s�EY͠�~�ĸ�s��c�����Q*�4e@�}��8s���7L\{��8��ۣ��$�Z�Ą�K&
[]�~i��;�+�����ӄ��yQ0~��N1wn�9s"T���҈3�0���'��� ���;ETAWi�;2 �h��~��q�e��o��o9Ommm��o��'��>��s�p�O��;,������|.��4Z_��Ϻ�ppv���"J�*���2�d[�J�/Ux��b�UU�W�����O6~yeu��O�e�sx��eQ!WZ]%�/�
�U(yU��!UT�E9Ni�O~N�G[�x&��|N2/g�8�����Q
���T�.�*Wײ��W�JW&Y�L�bO���O^i3�+_��E��'>� '���a��Ivzb������+���G�6KeV���Nu�����%��,}�x�Gc�S?��u+b�䓽��<��H�y�(i�Q���f}�+��}��זZ�c��]�J�E�g�51�Yg�n��.)9�=�A�]������Y��v�mf�k���'O�)��+k��>��*9�]m��b�.�0>��i��葤QY�-fۥf�4�s˸űi�P�SD~�r���ch@�?����O8��p]�`�j�E�s�{'UZ�q�v���g�I1Za|���5R�8��R�I����|ߥ�bi<���@ݤ玼�i�fk�8���6���<�3]�Sw[TVvŐ�'EW��زzc���G�&J==v�ܪ�ކ�ر�U�9�nm��폆ۣ� �R��p �OY8��>>���	��)�hn�4��/G�xKC�I3��G�Tؒ�Y���^"="�o�ԑh� c���w8�H���Z��'?i�._���.�q�	rM�f�6z֑ tp]����K�(�3p���J�c��)�;�¼b�S��h���!�n6	]��O�D�fCƌ@�ҧ<�� �]�1�ؓge/�.��$�fQW��b�T��cN���͏Y�_�/�!�\��8������g\��8�w������#ψ�S��d��D�q�k$�P�D��v��TjJꬎ�~ckT��'�9*�7쏖=0X��l������[���SΈ�O�SfƔ��G�Г�~�jw~V5蘉���c��H-�8Y�U�����ٹ;d{J��E<��4�(��?J	J�/��<���*�5��\�ށ����;x8��2w�
�ׯ_�3&�o߮�4�|�I�K�,�#FX�9"��*�����8�Ca�)�cՆ-�Seh��l]�c����U��`3b���떊'��
�"�"�@#'_�5�$4���9���I�6]ȧ�]`��o�ISV�����N��̏��^'�>#N9��8e��2mtL�2"&M'��IG��r'O��'O��3O��aSd���z��5�Hy�Z�@$L?�)�W�Mm۴�)��
bǶ�h���M�bǦ���.,��M�<0�Le3���WkW���o-Se���^[�(Dr�9s��q1��_nӃ�4G��o���g�/ʤ�Υ;~��\yE�89i�?��R�p�1��A��d�\}yjC4��ٳu$@�}�Ѹ���c�q�.�����ܽ������۶m��"�?����V�����3Ӻ�6	�♘yXH!�$�/k�Sb�E>��&��p%�[��,��C�@�u�O�����6%�n\�e��#�5kr|�n�+.��Qrt���R[2k���[(M�4�*�W^*�W��.���kc��q�e���O\W~�C1�̛��x�3���J���e��ŴH4��RG8#λ䂸��sb��kc箲hnlP�Do�p����x���c��U��k⑟>˟_�M��u�HF�b���@[Ӊ�d�ʌ,�����S2)$7�ʢ�yQn�����JτO
���ub�F����s!��!�G���ϧ�p��w��]�K�.��7�~z;-Z�	�ʕ+�?�i|��_�r�2�q��X�q�_�O���%�*����evMc�qK8՜t�G:v������ђ%�M~�H~s$�o`�2>IN�h� �1�yѴ�K��Ƙ9C�u�,�*�ZQGŞ�Rpʇ*���DoU�lO!�Ң�5�<f�>1Z+�I{�~mݭ�*�#��P��&��}��5sn<�#Ѱ�?sz�]#��y���QU5e1����s΍�'�ν�Ѿw�B/�w���H��*5�<y�X���S"���k�X� �tD��o,���ވ�Z�b�J�⡇�`�>�r8��Qׂ���R}n���:0��q�n����n�6z�eK���f>�#rX?Յ7uKJX�JC+�Z$��jqy|�{����+N:?� ��M��/e�b�s���Ƅ�!)
Q�HhA�s�S%V)κ�ju潱u�=q��g��?��k�e5�o)����l�Mp$L��f�؛�]jD���x��C�?��x��'�a��C�
w�D���Xt���8���(���x�GƠ��q�{n��m�����7�5O(-�-~fT�͊���<FN����Y��/FG���S>�F�@?�BЯ2�w��������5)�a�:�����Hs,���s������O<�h������j��H$�����΍G�Z-��	pڻ��L-�Uui6j�����\J;��W�r�I��Y��;���8^W=B,���Q�s:���&Z8!�\�c�s�%q���n�o|��x���ĵ�>3.x�Ǣ��Ƈ�t�uE!G��]t�n)	֣Ѥ�?�QWz �h����P���E3�_�5
�o^�:�Bar�)��3���ϝU�.�=V.�5E1y��X��3��_���"!�*;�[��'�.V��+�O�#μ(�tE��[%AO##l���kk�����şw���,�/�q��&�z{A��>�)_�q��7�7z�Ӿ�	h�_1|�3?��1	p:�7Wjd]�2�1���pMSR��/��̂���?ڗ ӽ䣰�DIk-���R��<H��z�.]w�|�3�/8&ͭ �%�G�{bֹ���o����+��x��o�5ן.F�hV���������𚝀.�W�e4��[s��pl+*��5�ٗ6�K������h��)e`���E1}�,�W��X?BVٲ�;�=�,z�룮�#.��E���S�q��1bHE?)�|kg�_�"�/6ϬD�J�KuME|��w��>���� ]�'k�_�_��ͯ����_�U����dK͕i����Rٕ�p�V��e��JZ(��#h�L�{�sb�ԓ&�)ި�R�,~�5D*1C#������+6��G�lj0��-^\��L:�Ё�q�o�	���_���փߎ+����1M4*��\2)z�Ѡ���N�C��6�й����ziN�p������5�t�|Ѱ��(~v狱��%�M��Ku�BS���_Sŵ��e�v�Q�+���ڣzbb$mX){��9c�j�do��y��Ue.[�=�,[*:�@D ���,%VU�������\kV�h8H�����V�����_�����]=�#����\>2� �{
ਗ਼ԉM���d. ������ὠ ��y���q�������R�^+���
���$�(�yqM��o��F�j�4I�<�{���<���[�f��Ӓ��ʿ���z\}]�Bv���lШ>Д�<Q�^�$V�D�R؍e�JW�Xq%��g�������o��Ͼ���Ҧ�I?� K(K̙RE���vwL9�6����څ���]Tя-\�N�Y8 �ZćF� <%u���!ZZԉړ��9�:XYiI��G��^s���� N�<o�w�W@�l:d��W�9�s��1��I܇�{E<����"��P�7i��;���p�3!|֪��O�e�M�LlLZ��q�������;{\\���E��e��z8��VL+���/,Y�~�_��u�f��m��T���WǥW_�ο$J�K���2��+����W]5#.��'��P�L۾�S��Yٮ�`j��G{�EIq�
�Ј��`+Jc��~$�j��N����<~��'b�?��ru,u�n�p<��7�"�g�?����8W���������϶]*���2,�N�&^��gQر%�������Ŋ7
�qՓ��X#�?)���]�JS8L9N ?�]-�-QQU�(�KǇ�N���o���6}�%�t���쪫���#Gưa��``�{x�}���q40�bJڌ���b�ȣ<��t9?
���d^�2�'���Y��kje�m�@�\i km1��ĳ�Z� JUn֑�1}$RZ�d��&3#Ǎ�R��B�@�d��L�d�ti��������ㅇ�����w�w~���'_����O��x��c��e�|����Ƌ�Q(J茐aa�A�=1��2-��TF#�T^L���ҨsR��M�ځ�1t�)Q5b�&�iP.�x�)S�ugGD�.󤭵#*ڷ��ɣ���
��xO�
ad@9�����]}}��g�Ə��3�-ԇ�=���³n�:�9 ���>���W�����������v�|~�w7��_�5��oķ��-o�<xE����I�9pU|�UÊ��F\�����$`Jo5���aƝ����y��v0G�y�-\�FTl�)��5~��w�U��U]Â_[SU5�d�P	�N�\(H�-vo�O��`�w�O�񇞈E�/�W��e�l����%���sO����x<��ǲ�D˾��R�xJC�F�:Kqg{L�>$j�͈n�d�t�)3bcw�/�g���U{���cb���e�I��0Fi�Η��SB�-�N��I�����F����<�-��z<�C'L�z�q��ǜ��8�pi���2Q@� .��"��[�X!�������=�C���'��͛����o���Â��6�̙یYA�X��hT'�T�(A�u,ڗ'���!+Mm���莐V2$���{%T���Q�HbP64�A\W�t��TK��t-=KBMG�S�����]�た�/=�\l۶'Z��D�HF�K���'�5t��+��c.�W�|(�7)N��6���{:����"�WE��1B�w�؅[�t������O=�?�h<����ƚ���=���mgal|sU�2�5F�q~T�M�q'��#O��kWjR)�סӴ�N����#�!Cb��11X�+#w���)��<� '���%ӧ>�)k��1'��ؘ8�� ��ɟ��l����⋝��\��L˺.��{6�R���p9	S��S�ї9�<HyK��Z�ڣ��A�l
R���'c���2�XW�F��t`��2�BH(_�^~������-]!M%:d�x�-�頴|����7^Y��
�5A�vו��*�����]�ʢu�u�M�Z\�t�W%Xl������<XQ&�	�(�'��zb���زiOlݺ7�l��6�=;��M^�L�!�Z��^z(.\�����q���c�+b��7T�����h���������Z�ݻ�#p������4|�6ɗ-v���M�'v{|������ٍ�/�<�`�TVV�(�-&�M�����S0>�g�#�����Uzf���1ֆJK���!pΣ���k4�Z��#cW�hr�-��,/�`����R$t��B�h@rT�hR)�]A7�v�?�n#l�ڭ����Pn�k]�|���x�� ��}����ѲkS�����.<��G$uF��*u�*�
��1<��`��#���Ӧ}��f�?���/.�~�x�?���wb��E>1�������&�
nӦ������W�F�\�)��d|�7!��p4زe�5*�:|�poءp>sʞ`���O�>�O��w8��\�i4ti�B�A\�|��<qr]��Pz�u:]sV�:�^��C�l��-��[haSú��L�����:m|V�����5`���y9>�X�%���aB(�%ۍ޺����9�~�]�S���:	I��bͦݱg��(��!o�(�,�h=��Q��#�ֈ��b�p&��=r���1���Q;����F��~��3��z��x:k�{�b���hh�k�.�#>a���.ndӧG�y��tq�����*��b�&�ԉ�w
~J*pێ?.n������q�6���/y��g�%���7�������˿�ڵk���p��U4����7��8'j\���� �����?u����۴~k���OZK-�D.M�����=&�,��$	�0B��I��b������di8����E�*{V� %�aY��$pشP�(�OJ�Ůnl�F�;�|>����A����I��gн��$Id����gh�v�9�c�̹Q^:8N9mt�HѨ�(ʡ�H3���(��䵼�BKN�$�u�Ac�P�;���]p���|Wd���QR�IjV�w� z�A<P������>�9�F����δW^y%^~�e�B��~��|Pv�Vo������zB�+�}��e��p���I0RJ1�[҅ܙܘ�Ι�s��� ��Ѹ�I��pl3�[�"��_��]���]8(���`�32ė7�:�ՠ�H ״�� ��+ң�҆t�$	��,�����ҖH�-��
���
f���,��=�o��Q�9m A���/���~��Ëb㋏�C��Թ�l�W3� ���ި�HR#���Q�'Ǩ�FGՐ���>	m�B5K�c����'A�P�V����;�;sP����/���~���n�!xjQ4���y+��v7I��"�F��L<�+���Jo�uƿ�B@vK��]Q�|q:��W���'�}��w�*6�rȠhP;�&�qzbsC���z_�}�A�oB*<9.L��g�K�wsT�Mj鬪�������w�k�;R�מ˟}$
Kب$ƫ�4mQ=-D�B��3��o<��,��83f_�^5ru2u�rB�bi��X��8����oZp{T��
c�e��s�����dj��9�Ί��^���#Ѵm����50:L��M;b��#b���QS�Mc��kL�^���
	�-�8�m=��X%�%1`@?�}�ۇ��7��箽���ܧղI�y����HP���+u0g$ܓDo�ϥ ^��� @�
��0-/랤hhn�M��j2�G���!�6�'Zd�����
✫΋����>%�p�c�ᨗp�rQ��ҹ�JJ=aC]�aD�p%��$�_�X��$W����9߀Kҙũ&ܐ�����%��ʒwӾ��KEQ�&�ʿ�;~q��x�'?����b=D���kc���QZY�F֩�~Ѽm�{ҴF+Z���G�����:�nȰ!�_��Nӱ���p��v��w�cА!q��Sd~����'oK�瓫_%<���w? ��\�l�Q͚����@���PT����d3Ѡ8�)�A6����nO���g���U�ƌ��w���4���SB+!+*�Y�I���I;��e��KN�С��ɚ�P׽��=�BiD��S�������8��qQ0��X|��5�Jg�BW�i�>�\y�p��.����uUq�MW��YK�ٕ�a��x��Pޗ�5�C��M��~P���(�%���E����c慗G�����CK���TG4��,s��_�4J�5�6v�.��on���ۤ���E��N�Lf��{i\��ۈ�����l��	����w�>��hhI������2Ee����:��
����o$�6)�R���I*�ԖE>� F��J°��1�[��|��4B�4r��¤Pbv��jl���]o>�Pt��*�\�b�w���s���Xu~=���|!���?��#b�ǽ�~ 
����G4�N(d5
{W��9`b�M+����C⊛��GO��vŗ*/�$��㖖�������ߤ��Z�^�?3�0����x��%q���QX:$
����Sw.���W���=yd�<Sxb��n���c�[;�m��lTH|�dN��������CSKg;n�����	z���58� nl��t�|�+�z��_����;��40�I� �B�� ���Lw鯴��m�O:�LK�Kq�8	9��F��Ƭ�8�2����<i�:D���ʲ���E&F >�}O{�����g�y�	P���+�O�������?�T�y|Ǐ^�����q�ܡ1�ߋݳ&6?{�P�� �H�b���E_�B�X���1������FiEU�uE�-	��(sYE���%������a9{��>~pwL���x�-1�~����(Z�T\�7�}?����&��ϝ[[�F�7�p��X�ʲ�Sަ��ػa���rY�ax'"����ދc�9�D��|\����O]��i '���Xsϛk��+����1����@ǁT��Q[��F��Y[��Y�MRtP>̃�▸�g���D���K6��4с SI���8I�����V�9!�*d���s��$�fjx��b���Ξ~Q�.3�NP��y{�f��L��#%o��;�/|-6��jt4n������Sc����a�ß,�g���q���q�'?ު��_|��س�(._��4�ܴb �EGA@�**��O��W^5�(��A��~���h�Ʈ��޷�u*�����8�=q�%3��fFT*������=��COkҷ+�(��%Q6`PW���D`�}Ѻ�ʫ������0۵D*���\�I/~?���W.T�	o��C�0o��!�	^R;��������_�d���ǟ��K��!4#G�t/����%,R��&�w.����-V��|{�It��mL/Uzw� C��)�yu�ќ� l6��8���1LaP�{�c���4b�䄡܉�W����Hy��n��
c���=n�l�IQV72Z�Z�9��ǀ�����[c��/ĘQ�1���b��1h��W_���i�Ւ�ѐ0@6B�]Q,�:|��8{ނ8s�91@���ʫ-�|�����[;��G�Ζ�S��U��,��}����%�*���(�����$���KTO��?n�7��0�4&O�C�Ŏ���ӶC�6C���ˢ3�O�6	%�#������Gq��>}j̝7/��:i�D�~�.o�9L�ùb�x��<x�:m�F���%"A�#�vi��S&��J��]�.n��Ƙu���qʌتΰ{ׁ/�ꀲ� ���+��.Ԥ &�i�����m���%\��$ \S8@kh���Տ�in�Ť����?'��h&���p��&Uo`��*�êc��cc�4e��qQ�N\'�.s[�{�;�<��u��&�֖Ƹ�FG����S98z�Yw����*st�4Rül�K.���/��'OS�jh�X��Û�3�Qc�s��om��O<$�a�/�R��4OZ���+6����X�����o��^��(��vꈘ0�X�Գ����y��7^�����5+5�jTM�ang�� s�
&)�c9:�)��'N2�SN9ł˦/���sX��7y�D�ۤ\Z�������}�	�Az���?w�u��J�:uJ����A�A���g������̀�#�v�(�y@�a��� ��	W1Bc���Z���W���b<�H+������P�կ�fS!�6C���z"C���թ��na)���DIG�<qp�=ғ@�'��`���f�֯(���vQ|������������">��ĵ7�+�:kf�O�uHhT/h9��<�-� ���uǊ%/J��e�5�+MIm��55ݝ���щ! �5@�@�c��ĲM���b�ֆX�j_�X�.����3;=�;���x?DS/P�q B�m��xqѢX��?J:l�x	���r��o0
OBtd�U�.���z������&l�8��ӥ�b��M֖G3G���n4~�+� Y�:	�s)�!���It��t�f��@mm*�A��x_[�;���=Ѹ}��]��.�y�F�e�,�{�Q��[P��M�ld&#��jm�I8��E$�"�3x
��һ�:���#���~%1��0TtEmyw��HH;4l�鱓m�������
��I�;�${��ͱm��(��+"��/~�+z �|H?u��]P�k�7l_L��<���Fݔ�c%�z�e����+�F����0�xsE����=f�F��X�f���) ��m���$�W_��ytdL����۷�p�􏪪�(Ӱ�ɛ`�p�@t�J��zMb��L����\0Eh��([ ����p��2���N�ΐ��M�.I_�x]<��=Ѱ��kS�a�b� :���-�@�a�CY>���.Jd��*�!A�a���?\�I\G��&�����-����Vс�e��:��U~��N����K�}^6�V�Q�*�ɟ��k�JQ�q�����؂�rb�����c1}|}̙;>&��7l�`/����e��q�'��N ��I�5�^3gΌe˗ų�<kE��zw>�y�غu�1{CGuu�{���C��!��@�+_�P�-�M�f�ZX� �m��f�$�0Ho�(8}�$c��^ol�n?���O�P�IB�߬�z�5N�����D����Kk��{�mk
u����jKs�Z�~o�
L�Y�eVh��',�:��ް�]�ui�|h��'<>vZBA
N��,H�Ѭ2^}����c������
z=�7Q����]V[�ۇ���{��Ǻ�k��a����I��]'��&e&�#@�N�y�Go�yú1|�&��M�; ӟ�M�رc�B!��`�G ��o���?�Oi�m�~�z1�'n���#��о�Sٕ�h�8��Ò�cQҴ�	F�
Q/۷�K�^ܔ�.�~���@�Yx�) ��P�3(���֞x��Mq���҅?��Iڕ�C�$���x�R�kI��G��*�:�Ã�o�HP٪ȟ�]U�%cPf/��tJOW��:}����Ԯ�?o1/}uY���S�Ѽ/+�t��.,���TQ�<�u.a'O�&R�b�eWEM@������1|tM���*W�]���>D�C@h�H�!���{�͊�;`�|@oW�'�vő �DȷK�7o��?�л�:�;�AvpYyy���x��'|0�Ѡ�P�k}z�@YI��߂��X�t�P����3���i��3�
�o���kM��׆-�q���~��b�'���5JT7ڍ�{�:Y��:�s�W"����_�q���:��9��>	&��m�bCq��E�gr)k��x�������-�'~��h�-Ӂ�t
JR����\rY),�^/�2��(iUMQ�[�-^y��X�ȳ������.��_SU�5~�Q�H�/��މ�6�� �x<V�\�����<�mm�M8�����mӦM������iR��ܣ���r;�ٷ��4���̑�=�<���^���V�i�E�&U�t&&[�\�D��[�Ӑ��hm��q��h|K�����G���R�0"��ݨ@OV4�:�(N=krL�3;����Eu���i��b&&@eMY<�ěq߿�C�1�4n��ߍ��#�e%J�&Vyؼ�T����\\*a�9'��!M>k��=[w�C�=o���Xxs��Q�C7��S=��K�@�zZ;�F�B�\U�г uʣ��0v�5I�#�q���f~��1I���Kc�m�r�y�"�Օnx�[ʀ�9��2I�����=�� #�ذo�x똓���o䂣�J�)R[������ol�vi�TA	��p�31b��W$�#��jX��=(<�6�+]N�aw:Va\���?�R����`�&�u�$�l���-�I���}#�M���C�[�!���<|���_��O.��}����f�P�hP}�R8�8�\�K��N�w6���er�~k�M͍�O�i��oƲǶ͚0�����UM5d�L����M0B�/���Wڼ������:5� N�/ ԘA%%�q���F݈�s��2�N(�0J�� ��4x`\t�EQQ!e�w/��o۾��+�F���=~|�C��W�����$AE(!Kg�}�@
����,�B�&<c4��,gT=lҘY�89�<��,�w{p�$���&��'t��1h`u1(��5��k2;8��?�!�ַc֔���+�k&�E�����<�`�L�����DkkK�5쎦��ؾs�&So���c׎�����iJ����PI&>M�-\�*JK]�ڸ+�G���]�h�
����V�4n�9�x�BRzx�yKiYA|����]7Jq��S��A���O���"��SA�r�g[�_'������~񟥁[�3�d�Q<����%�����ӆ貲r�kB%�{%+�G�o�U�rL2�"����<��t�7ُ*��8�.�4>�De����8j�*�z@ml����^���ٗ��U�T~�M+�pq+�K���[Z�Mu����%�MQ��惨}4����R�9�G]L�HB,Z��j�M�k�I��$o򓄊�Nm-2�:Z��P�Ҕ\��2�_*�7�E\�)�;`�A�������^P��,�+��sR�#�ܮ�U@^����^���G���]���F��VR\\"�W~ds���x'���m�������UI���D:SJ������(@���f-�7��I��')�����Mf%ز��G�ւ<�!��;+���2~�&������S�`�(T�>����!g�۹uuW�[�{J7y��i<=p��6{o��D� #%R��(�?�i����!�S����
X��)��I��qx�L^���`����m������j�t4�Q<B�����}e�&��4Xؿ�)x�hn#O��'iL�}!�_� [�t�9QV^&-v�,t\�g�S#�zE��"��E�rEp��it���ApᄫJ㼾��E�H�F���M���UZ� J�*T�H��[��|�QgT�p�Z)-�tM���x�͛���)�ps���ɗdF�I��ȳ���;ڤ�ۛ�@��4��
:�Q�P�������7��B��<�ł�D>v��۷�0^F
js\ ?U��c\�sްac���>**9d��`�$8�3M��U��@l��5kV����
�uD!&UQc������t��lT	+B-@V!�x�f���T&��/2���&0_�
���xx�LP�|�C��Ԡ����4�	�^�>��q��q�&-��D)i���)[i��*�w��$._ߵ ���(J02��ʁ��G�R���V�Ú�,̄K�Y���ը�Wi�/(���סI\_�¡�<��͸S8gR��C7_���&�pF �=о�O���^��A�-yyI���[e٫�[���ĥ+Kh�/8?���Z� �=����D����c��S}�.�s�W��!F���Ԇ&(پ��*�BJ���4H~o���MĦ΄�㓦 � ?���@(�Y� �8���O�}t��F�!�S�� �ҀL���j&j��h!ҳ���d&�N9p٭�ȍ��q��A�9�����e:�$s~2
rҪ#32��j�,��8~RoJ��ם_��Ǩ�/�2)����0��s�SO=%{b�L���ϕ��� ��qB�o��1q���Q�i=�8x�3�X��j}D��a���\q1mIpT��B #~���ٞ�-	IcT)�y-��#��,`Y��;Ҥ�$$�S��LB�A��t��E!A�^����W��lH�"�+"��˞9�>�N�%@0��S�"��'8��C��.8~�J��4C����p����@�;G���<�j���U��c.��\��>�����K.�~_��L�C�E����{�.1��!��+�ga�'�Q�@S���<���e�Yp{bda����;�Ɩ�L �k��.��<�%���4*],��|����S]w�B�1�+�s>F&���C�NNX�;,�Q��:���_BH����{�g9�ӆ;��J�wS�X	���޲y�MK41B�|��ȿ������;�3�HB�P?F����ω�Æ�@_��}����Ң����m_1%�D� O����\Z� ��4�骡�'cƑ�҃��V�'>R�{�DR��L%�!��H '�%�Y��њ�0�����$Q�fn��q��C%��5py����JY��Tu8|p��qf�9un��97ƝvNL8}nL<s^L�� &��Y��2�1�Rݨ��(r�r��m/X3���M��֤�nx�\&0��a	aJ�� �>xР(���Qfl���sD)/�2���o��wC !^�|��V,��ʣM���/��>N��(8�$o�ѰdF�y֠�U�@9�2�ȷ�E��8�o�#!��w�C8RLJ���M"?�`kc:���M���y�[��%��^m�-͚�񲥈N�Ң�0�D�������8������0Y$AYIA�?oJ��ɛ��@���7ƭ|���-�?rc���7��W�&6�du�.B��)\V�'w��&˔&��d2"��ҝ���6���;�W��N���#�4�yg@=�VR^�_)��(��~������{+{0p��k��//~�G������<�J�W�Z'i���K/y�Z��v8༄Uk�D{c�p-M<���&�Ĕ�:�E���B���U�0Oh��Z�� -\ŧ2ɨ��l���#�N�S��g��ϘSϘ3�8;��5+&�:+F�4#��F	g?iA����;;�,�|���46v2�m����4�;Ad0�N�ߖ;��11r�T�T�g�O2�y5=[�v_l~�YDm��co�.5ɥpg/��&�^ć�?��(�����?8U��s�iS�Q;��q�1gG�=Z&g��R˖.�J�.ϑ�ƎS�L黌�!���f�#A���E�L�4њ�!��%7e��:[l�p8 OMϞ����c�8��\?~ş�|U����L���`qEN�Z<�(�97TUǻaG�:�):y�n�Q1��SbҔӢ���A#�%@��QHݝ=Ҍ<�.�w����ZZڢ��=6n��o�7^[ۖ�rk���v��e����la�BR����o����ύ�_-���é��H�DYmy��ѝ��7�Z�:�y̰/���d`���3��=��wI��Z:��-�CL$�!$�E
 ��[Z�c�\oolJ����rϐ?f�X���bٻg_�����ԫCJD���K~��x�q�u�д	���!��ø��0�޻y�fk5*M���/�9k���u8��k�IM����;Ę���+�����ʙ�֦H�%����B���BqI����߀�1g������Ƽ�/�	��F�A̐;���U��ow��Fssk�67G��
	ڠ��qʴ�q�sc��Ih�Yh�7��7����{;��L�XwI��'J����c�T��gv�x�`��A�42 ~��+N$�	�eGn�/$�rL���tq�������+��Qt<3`C�]_�a�k��|�K�5z/��˖�X���F��s(�<<����	�&��^a?��;b�/z�I^�#�+���yz�a�Y�]>�b�@���'T|�a�Џ�ҹ������Q`&���Vڜ��ra�L��U&aTyuuuq�uWǔ3��Rd��[�e�:�)����,�*w9h6�	� �ZU[�^���ۿ��­1r�9���~�FјH��F:[�=�/�JĶ��0.��8��w)	��c���$啥��gw�S���QZX/D{��%�8�C�(�§�g�lrV2����g�4�fز�o{�E1{�5	�k�]�z�{֦ݡ�Ό9�2T�#�RfN����g.� �7!�: �7��o��{�}���~�$�iB�D��8�YDl�c�j�脪�'M$�6��J.�(�����at��*-�짞��7�ԙ�ejB&��ࠒt��|���0^���5���H�M��	�&����űxŞ�����7ƻ~����kR<����y�+�[�$��hE��#@FМ�"�5%�q�5s��o��"M�[��[���IWZQ�?�;���磴`��:�~�(�+	�w)fj����o�x/�Ә
�wħM�}⥕ �B�����~�OuK���B�K�I����O���*�*C������W��v� �:��w~?���"ܢY}`?1�B��r�e���?�%�����$SqǊ6ET��>c� ߋ '�Z"�Ͽ`^\|����C�͋���8��+C˛�e-[x����\]J�ϤGM,��!DU���7��7_��e��?�T�ya���%���Oc�ʅQ\������L� q�Hе\���ώY�GeT�cq4���a��K��V��O�'��s��{��X4f�� �2��e��x-��:Z:$�i3�p<��V��je�u|��|�{>���Jm� ���ƈҭы�/<����8 ��h��L^�`w���_1���߈;~�p�k�nm˘�G�Xz��"�S`0!�u_�H��y�� ���`U�Fc�'b��q�-�E�a���X	Q~	q	+a��%����̼�Y\�Nt��PȺm�ٺe��������}!F�����'c��y�ݱqwG<��gc��OH��B`��As��i�GցxN̼�ݢ[&$)����i��ڊ��3{eB����t|�/��ēǨɫurqǋ�l��MoS[���O�r{�_��R�ʿ���f�2���-((񖭰~� ��r o*WF�F}���yC�2Y�zߍ'`V��/>k��� ۏ=�".�����؝FO򎱌QG�������c�LދBh�f5��t�1R,�����Ó2	�׬A�"�r\PHV%�ʔ&+�UcH�iX�R�x����is/���/��((��d&��a�KT��;5�gy��\�Rr�D1T
Dh��uIyI��Z��_��Ek�����1e��Kv�Ʀ=�胋b��=�ޔ��
�!�\�!��//��̘u�{U��l�B���ˊHui<�bC<���J�����Y���7j���.��k����@G�	S�s���;�D�S�WC����b��h����@Z�'����&��j�ի�myƙg�X�-[�ƒ�1��Ul֓20���Lݫ��*����l��4�]�É�f�}���+v����B�O7��]������Vqn,����yt�Dnz5&� ,��$JSu�PH�pR�@+�s�zg��< FN��� ��� �@��z�T��)\Z��t#�[���9��H�J0.Ũ�[�/o��G֕ł��Ą9I�Y�{�A�M�vz��Ц���ED�ǄExS�SQT���l{�K�k��uڔ'2.PC��5#0yz���i�$�FN��W�Fr���9L��Yj��ګ}Ĝ�g�!+]|a�w޼;vl\|��q6q�Ї�sPe�yG�q=H���h0�ڴ���W\y��.���v�Yg�U�\s�;׻ӎ
�}�Crͱ\(�{E�.�@���&���G�\��;'��P�Iq�!?����â'?�m���=X���nW��pii�RV'd6�B��W$��bc�/IT��bR	~������q�usc�+���_
T���D+����s��$�E�.�U��:�:���.���ǎj*�a�>@Y�&\A^қ����`�jw4�Gp�4x��� ��[1j��v����z���>�g�>S�sCW��nJ�_@9� �
b�i�y������ӟ�5jT��{�1;�����:$;�PQ9s�����i1��+-ɶB?�B�����WZE�Jc� <=Q.�`��QQ��x�8hX��w����恇wh�����=;��7^���,���_����Q�Q���,�ɓ7?}C���L�*����;����;'&-xWtD?۽�C��^:��С����׍����&քȢ�`�r~��x޽ȿI�M��P��	�i�J���>{MA�&(�S����%N�gu�'���ѯ_�1bx444�� �㑙��X�*c���vT�|x��}� Q���׿�:~�3ӎ5�4ST�^p/��$���T�Xm)H4�!�0Ѷ��8��M0��Z	`�Я�6�w����E�@�$�+���^}%��[ߍo�ӿ������׿����������g��J���a	��(/���b���9�|&��H�:|Ag����b���^�X�Bɭ���v�]�������l/�]Jc�"���^�=����E�;6	x�N��aXX�:��V!|�2	ѡv� زiK<��C~2���e;�*Oq���*���2�<��Cz��^6�A��8F�ǿ��mT;� <��@����K�pӚ�(5�F�K��kB�D>�~]�� �y~�Y@������a��^:NO��G�B��{�����xc�Ruҽ�صK��:b���X�����w�{���x��G$�L�Ri��I��,�����i��f�*���%.�vv�=�B5\���<^b��$Y:�����+��Npr�:����ũ�\ə��Q+���xy,��S?�/W΄'�M,�CB.�P���x�y�hܸ�ɞ���iӧDKS�ϐ�ׯ�O���櫝�F��<�X.���~�c��e����On�c�$�}�[��e�J�M���0���,�'<�Bo����^�J����)��bn�!��rI���!䫮,�ں�y�2A�V�¢�X�tu,z�hmn���Ci:w%� Vį�ֈ�o쌟|�g��?���="_u���p9�(��I�Eg��%���y��ug)>gJ&���+�� ��� �������p����a��?��4&�o!�)8w9�8��3Y>����H�`�������?�Kd���l]�	��+h���\�b��q�d�h :x�pjl�.\ z����0/��8}�,���[o�4rG��G>�޶q�F��,\ʎ0��LG�r͕s���\�LZ{��2�AՈ�;9�x��k�7~��c�P/mh�1�&t!껈��6��+Ͻ=m��(Q5i����gQ��=�:��ߎ��}���!E�S7��cT��)��ɣjc��zԩ�'�L��x��*Γ���R"���!�D� ڵ#1��tdIB�H[h��ݦ��	z5u�5��euPı��!�+�^�/�RGe=���65�[�lY,^��������Q!F{���vl�:;��d�~���[o�����Z���b��o��'�x�n!:r�\Z�k�m��ͧy?����<�Q�!	�����X�R!ys��bOVYB �F1bPL�uZ�TT[�!��q=1Ԭ���G���$A1r#����U��K:����;~p��2#:�\�:i�ZB�(�➯�/J��u��EwӶ()���?R�{��D�pH9Vʫ$�%��n��gU^��g�MN�O�c\t��>�A0�'|�zB�+�I	�q��i�F�öESs�O*Ŗmn>�������w���߰���0o#�����,�u��5��wX<}\Sc�˝q��1y�d+
Cڻ�*g�	038��ч�G~Ļ���δ���x�'�Ei(pP
�Áb��,��"�rR�M _o����42( v�B*6�[e��̈́�6��\l���X�ֶ�j��� .��W��}�F1J���R�R�����x��cŢ{��J4(�H=��@4���6.��Y����~�l��iY8=��]��f�t��
&^���HZ� �GR9��#�Pp�4�
������S:�It:����^��Ǿl�������2(����$��c����pnА����<��$��[���7��I�
��{13ܾ���&.8�` ���q���_<��f��>Z)�cr���uFk܌�i?0G
I��h�E�%G�D�2���/��o_�}ִ���DYe]�3����j���x]j1�������g���Ӕk3�hr.�.����Y(�!Eg�ʈw�o~�8���,���N�.��T������*CG;��⎻^���a\4D̽�f�����՞��ZH��J+�ㅷ���/��F�͚#'��|b]�z;W�TL��]4��\����fb�_pKe����w��ψ=&$�Y�$��Î�A9��:����S��n��Ih���!�Z�������_h(j��i &Z~��y3�B@�MڳD���jSYi�(��B�����3O�W�z{����6f�һ��D�h�\Iy��ۏ��ߩ�j��N�+PK��|��G	�k�o��QVS�Χ	cEW\z�9q�9WDA��Uh�b�m�nF*�y��D��j�����ڳ6ι�Ru��	�T@e��ElQYa,^S�~�o$�DCZN�\���sD�HB�:�ыc��jmT0uT�\�I}Q:��OQ*ܝ�?�����O���C�����!�N�*�wn��/|)ZZ9�Gcn�Y�򃀈���  j��z �ՙ���	�O�*r��1��$ ը�s��;=������ػv�:=���@��a��UJ�XU��3��K�<�ok/��vDYq[6\���4s�4e��z	k�R�1t�`�VK�Eai����3�,h_���ě�S�W|",M�ERFh��xCy���_oT�m`9w]ӽ�X��D.��: Ι{�����x��(.}�.]
'�8���!칉z�f"��(���z��;�����������p�،�.P#0�cm�)[��JC�c@~�5D��QQn����J�����u�pT�����	�)Wy���?x"V=�C	9���L4�ˍ���D��Ժ�Q�����2��S��3��4οxvL?��(.$b;�M���GtT*�P�9����V?�f3S*�o1�n�;��x}a���>����*$�Q��?^r������'�m���f�$��)���t�Nx�I�"�@^}��8����@G :'�b���˛?�'��&fY���c�8�..��R�-�
��}��o?�w>e�8d�0��\��g��UTV��=1��+~��˱��A60>'dLW%i@���F,��	��ҵ�N��=as9.1��ƙ>ix��DU���[��J5�Z�tJ#Wď�x.�x��2-���	E`�#�he$�,?$&�*�*�H�z	pe����sN�4C�ƅWʜ8���*����HI�)���,rm�@�c�݃�S(a���ަ"��卅q��?'�{�4't��.��&�t ���闳�`��u�O�Uz��j�$�3�D1O���L��S_8(���5v����xT�r+�T��>c���jW��]Ҭd8����=7�'�͛��;�[�f�<���#:�C �Kv���b��ϊsΝ���2m��I�����\��@8 �C�/&���&d��#�h��Χ����Or�ى֕�E���3�>����ʚ*kb�c�7^0a�� e��7М�HX��n���y*6�񨴎�5�	YJ�����8=y���`�$U27\W��R��[�������͉��YP���g����o2#�2)��>����Y6����/�8>pۭ>͉��U��Fĵ�_���q���]��p�J�XIڻw�ir; n��������G���}��<�[殿���Їn�k��&gGD7��Le[��"�,�ZJ�в6�uCهP��$w�dR=I
g�߮�[S��T�|A[��#a��)�(r�U��"6�#��E^p��=�@��sշ��%2D�RM��c�N�koO���b�[���JXI��٩���y�JB������Fݺ��T.�X@��ip��z�H� �)��вI S]p$H�)9n-���u#a�?i�u�砌�i^|�q�Yg�뮄Q{�,X�-�pb>�Cf��ɽ�W���a^�c��	�A*�X���W�.��>�g���~b�k���n��|Hmb�[����h|���뷪;`�-���DMz�YKKg�o��!�D��=���tBi� �7d� i�Z�Ns�FИ5��ʝ��AՕ�X�I�]`!�֤�0��鎻���ز�)�~�;-�g�`��`U�$XB�#2g� ��n5"j�U�$t*QI��\3��v�h�h�S���J9��Й�Xp��〜W|��aOq�<|�+��q�셼p�|D �p����{μ!���7z(��z�k�G6�H�T&��\��v3m���@t�^r���=�2��*���!4	S�reii툽��81�H�*�aV������G������(�!�����"u��"./�cxrʟ�'��o���<�\�X����ݸ�%�f�O&����8*?��ɏ�5��B���R �N���6�9?!�rśG���l)��;4����ο�$�x��GBs-�<�Ʋ7�ǟ����7|�	�_)� ���K��������"f�
1#��L6e�ٵۂ}4�`����J1�F��0-������4�	��@��� �-yُ�G��^�vN�'�e	�V3�~����ʤ��Ʋ �+�K{�3~��_�=I3%I�;� -�j��X��3Ѹc�5���%�K�`�ө��&�T$�':5�)��"����i���0��G��H���m�� ݔ�}�c�g��q ��r�|�rO�&u��9b�F���#L��܀�����n��Y�� O��8T�%0�C��b�8��M�1Ne1s��S��|�XK���JX��_�N�ՠ`�"�T�d�wJ��龽�^Aj*���@�*�����Jb���T��(ByH�9�4Q* �f���{)NW�BK&��p�R��W�(�-��?x_4�]#���H�
��8	"bk�XaɺJ���\���
n���@	���=� C	=�����Kg2��'�)�<�J�K.D��_���w���A����&��L�(�g7���������\V��9S�\z�����T��m˫D�}��V����|cǏu�6��襵c�7���x�fƫ\N�9�}b��͎�T���&��L҈�D�Ҏ_Z���g8ܴyW���E%���"�)�
K�9���
���
 O�r3P̴_���W�w�S��b����6oT�=���x���(l��l(;X�a"Gu
��G��^�T����.���)�ef�YL�I�'��K���v��rs�Y&2/�� ���wʔ��B�����ؐ�C,�����I~hk���sȣ��V��-�.��9r^�ٻ���E�^�&�(��g�yƄ�| �-������ML��U4��K,�O<u&��!��v��	��� �445Ǿ];����-�ow����ƛ��fM�J�zt��8����3�Fy�C(���T�����/���zF���m����J�����K�%��F-�ե�P#hRRS��n�Y��Ο��E��h�D9ʔ�p�OAB�&�>rI��Ju��!=vN
u�c8p765�2�ʏ=�x<��S +@Կ�r�*?�c.B�����;-�;+�N?��și�dl�M�����<���x�_���<��L߹�,�����x��%���1=�3��D:�+Ĥ�-���|<� �Ӑ��u
�D\Hn.� 4򕈱�N�O��}0S�
�t�!��**���{ֽ��ӝE(DWЃ�F�,� ���Y�u[TT�Gqy�ڮHO�Y�҄΂-�P��u�շ^'ϽJ��l6un)�iU�/��S�*���Bt5.դXI�@Cz(!��Ӭ<�e��0p��&�|Y��a��9�ץS%	Ma~�@W�5ώ]�).�:2�������Zn~����yI�H�������>g�=��n����}%��&fH���ґ�oT^V�,&F���x�ٗ���)Zx�$f4~�cZ��xb$�<+���є�����wb�@q0f8���e�L:4�1��K��-�/��_��(Kq��<A�V�F977�(ok�W�G��&F�T�ǁa2�B�r�D��9�<.�1f�<5tz��ڧ[���4:y��7wWķ�������]q��d&���q�x^'�<���c,��J	Y1��,p���jD7�"�.��}�cN��x���@Q��"��h����+�'�c8P��͊Mҷ��rPi�������{��:[�҂>D�򩌆7	�s%D�0*�Y8L6�
�p*��-3Nh�ǭ��eu	E�iB���P�p/�����X�ٟn�V�� �����Y�,�G��X�Z���Lxh�{"��h��9Hk��8�1h�d��*+�g�hg����%A�����o�]�kNg	*{�y�a�����{~�D�3����&/�B�1���O���8�1�>�/>������A��{��A|�����[�4Kߥ�����4.'�`JX{�YR�@7�쫂{{�� �,�NG�I�ߋI݈@��?���-V;��b4l�4ʣ�F�':ڢL\�fE��x��<�� �t����؏4�dʕFIY��(��nG�(�K�+��kW�ilB�gk��x�$t�i�x$!N��|t���V�=_�ڗ��� c~�*x��w]�7_L�@� �����pA����p���|�����׌SP.��˖.����W�G)��*�ԃw�]<���6H�R�A��hx�!������ՀjL7���|p��szMW�FK��K!M¬�JO�L�N�mfc�L�;uM��O~	�d*��7&f7;��� n��x�$?��	q^C����3�Q����7mHӧ20t�=;gGBp�zy�-ǩr�Zڣ��	��:8����^a�c �Iww\q��8�܋��9@1[!��/�/�_L#L�옣�؍�i>�90�۰1�泟�);�vq`�͛��R�8�Bǳ\[��>�j&�-
|j6�:�ޖ�	oI���}��ꄩR	R���t�+8�4��$l�EC�@�h4{T%q^ew�Ʉ��W��@��֞D7�o����c�˫��^�T/�QDyd��(��LR��L	 ;	�Qg����/�)��e�U�*�W˓�?�i�7ʪ�P�k�<�f�+�|n����+/��Q��|��;���ԠNͲWUM�������ş�e+�식ei��� �q˭��`���U�$X=�mv�gx���?�=��Vܙg�Bh�������3�����h��n�g�&�+�HьCD5��/�!)Į��?44a�T(	q)@���b]Ɇ*cR��L�&�g��!�i	B�Y���X+B��&ۙ<�,�Kw W��O<���_&CRh��z�&y-�����wN��?�G^��� �')�F䔦K���ώ����@<΁��,���^X�6-��Ϙ��L�l۶m������\	���v�]��G&�  `<m���4���ٮ��*O�����>��8m�i�+BG�d������R����r�K��D��M��U6��*?�mͭr-����kS\�&V�r���ڸW����՟�^Nq�&�p�Nl�
n]ە��M�[ۄ��y9�S��G����{��D�_?j��&x��Hڧ��o`��K�J���7N�Dk�6KO֜��C�r�1�Ь\�K���p&AI������'m��@Z��k^�7]��xP[��8�#9�O�4���w�!L�N�7n\����G��;８u�i^�U���ʝG����G�C���WtǏ�O���Ɗ7W�l����nnN�����81F4|��:Tx2�ΘX�dR:��͘4��ni��+��˯R@YEyԍ�����Lt��8I�}ڜsc�I�G��S#��{g[ʛ!sy9.�hd���MD#@ŶY��Ht1,N={^�{�Uq��+�k\~��q��7��w�7N��t�h���L#+/���	�I �~��c�%��x�|\,�,��$9�d��K8��\�I���_���x_8#&���!;Q��+����:�r���׾6�dB�0�"��6}�����>O?�t�w�}���ۿ�3���+_�qAG*PVP�=�r�G+JK&��Rc�$ ���
�&7��A����=�޴i���;��Č$8�{�Uˏ�8*�]~e�0-*�*�T��*�����@tJsj����;+��S�pe�db��|��w"�a�4g�1!.|��c�i�cYp�����˴(Qy"�Cu{}G��?���O�De�3�� ��;	�li]�Pr�dT�a����B��S��s��#�sr���O��v��/=7Jk�pT�y�!��R>n���ϒ�2��|�M����x�7=�;�w����]	d�<s�/uީ
�=*n��-�q��x�������F�$4���{�'�1�ֽ{��,��#����#)f��F�lr�J�p���T��@+�Ƌ4�&��麘{��1q��9|�����ڨ�����-�?F�W^17.���(�a�f�j�raZ�#ڠ��i_�꒸��kc�s�P�тb�^��`&0�����(������Q1�4��8�}X��a�Y���i�(����b$���
��	���3��v���W!j���cC����♧�����5�̞6q��M7�/���p^Y�G��yvx��1[p_�,�5�e�v�暫=$������!�K�M&�&�(@�^GՌ����W"��y0�Z�0h�/�I��'A\�z����]a�o�2=	��e��'�c�O�n1�/����A�c���:�$��1V�\;t�*�n.�)%�)����Ҍj��c�ǐ�3es��X����mRw�rM��fٌUE]1t�D��&�p��Px�}�4�CUjG��%���}����E��<]�M���/�r|�uW�L�0��N���/8�|s��M�����rp8b��=�_�[��	�_�<
�Eg�a�|�S���|�#��,kp��������O=�(��F6wz�<P��H�e��jt<������ׯ'!J�Vb����@$�'L��* ���{	AMM�?N��~Y�S��>�=��P�{5�J������HH����rŇ@%��Z��H_%�cH�zݷ��C��&��,[D�Ҟ9N���Jw:�i8���>�����-G�DS�%��| �ȟiSb�=g�b��e�'B��q<� �JhY�`� ˞qܠ�=i�8��8���ě����JT�2
�i�}��w�uw<�����ϸ�p8ۏ~���ɝ?��_{-�#��)��@�	���r��<��x2M#-L�rm�M�~��m�xR������?���)Iq�i�uXja-�ɖ3a��v��/)�*+����*�!�/o�}�ם;�wH�P��"u:��'SH)a�0����(��u����RXQ��}��[ U��c�O$)�L	�Yޛ.�U��؃7�f��9�ǌ�y���/�K�^��۶;��h�>�X��i�b���^���C�����;���V2�8&T�=��5	N��N)��d3��3�����U*p8 ���9�x~I�{�9#N�g�&�8�Io�ꞆM��Fc��w<
ȇ"?����!M�]�%J�T鯺rn\x�mQXZ�Ǽ/����T
K�VSW �.(/�����o?�����b�Va���Kh N~�htт	q�}.�:��ҡ"�ˠ:��Y�v�a�tEEMe���Ƹ���Rv�v�S�7帎�P�I5	���k캋��<��p!2��U�H�
��.8S�\�[0�$�?@�?K��@�e(6ٰ��j���tMN�͊?,�Bnz�M1w�x��������+��RUIO}<��b	0�b��z	���I�6Z^9���˄�M�<��Șp([�P��Q#y{�W��x[U����zcO��*����L���`d++�������=�<�}5nsV~*��\�[W����;����������]#{Z�U���������i�7D���q�������(����eU�P��(�-�r�r]�ƌ�T{x,G
"��$�.td�m:��0�L��wZ�~ΥN�Bƥ���~� �̓8����m���\��ãb�$ �=J�0�r3�W"��o_�l<�̢�o�K�-&L������|�Si�������M#��_�G~:e�=�RGQ���W��v1w����j5f�����_�q�
YTZ{����<K��ڛ�	�Qf~~�� ��:�9#��w��9 iu	����+�T��I���I������~���7��N�.��<&���U&,�r-܂#�f~e�p'�=tE�PiM�v�Kϝ���-�� ��(��0�����0����$�uu�����:�Z{�P5VF0�zIp`�n�4��*5*CNm��C���	��)
AI�61�Lt��)SF�]��4&�rG�Ȑp'`���Z^mk��DH�I�\�E@('9�76�d�-�J��(�
c��Nuu�T~���z�cז=��2�H+��'�1Lahoo��Q�2�����K:��N���~;�AJ�/��`#�XV�u��j��=���Ƌǋ��`���k_�Z�ٻG�gP�\��'IFE-�8˟Rк;}nq�o����*iX��pz���-�y�h	/�Q���
�S(��r�m�8�mᑣS��Θ5.��[����5�p�GG_��2�	1� �]Z^+����wb���_�#~�v���#]�BT^�4��!��;�{1h�ݧ��c[�Ge0a��hv��A��)�o���c�[���� ���շ�������M�uo<���My�tF��<����@��(tɼS��nuބ!���@m�v��lD���{�F��u'�%j���4��<N������>�E�N�K����h
f�<�7��F�fu&v00g�@�jJ�$�Kb��z�G��n|qK���ʟ�O���*���D�Y(�	�.��ȟ�U� J8f�pT�������.���薉�&��DC��$v�T\����~�0��F{�V㱩@}%�P�
`2�6�:�5�h����q��?��DQ%�~ų%+�čɰ���s�^�~�z�p��ӱ]�]Y�OI���y�u�J٣�U6�Eg�D(�~�:��'o��C��Ӽs�Ŷ�θT�U\����G �>�0@���F��:'�D�%�J��Fs/��q�Hx�=��7>��8k�Y8�|��h �G%�7/��s�����s��:�K�ǒ�_>�JpT6�cϾ{%���ބs(����}.� w���V���,��85c���Дm��,��1v��8��1��Q1`�F+^6�z�&u���xUu{���c�֍B!R���r�˥Q���aF˲�R��'���'�u#F������
�8l{��X�������l�� ������4:���sT�^
9�>��}}���':���1(rɹ��?c�bR��8y���Sf��D|N Y�1s�7�pp��]�b��%~�!�s4��Q�n���	0�b��W]�\vi�ڹ+������x�{n��sf�ʕ+c��/Ċ7ߒ�:���$�M�����>�e4 �0�JL(�F&�G��i9�d�f�m��x�{~' ������nCK[JG8tAsUmU��.+-*wF�&p����-��ũD����0m޴�z"�)��tO=��ޛ/�gV!��zC{ҕ�+Y���;������_��!J�����x�{�6��� +q>�7z��Z.<��4j�Ï�ȑ#}��	�ի�;���G�/�Џ��N9��Χ=���Y��hi�|Ի�zkpd��Dc�]�ƕA���s��R�y�Y����P&@�`ڔ{1Sv����|�� �O�pf�|�T0�f��P)��@8ɑ]�l���a�޹'6���V����W�F1~����}�hٻS�HC��YUF���-m��)���A�;{��b\g�5������KL��0�7���Y¢��=�5'�;�$��ӣ%q96����0����J5������Oy��i��خS��S!s�!��� �uͪ�~=�aG#���p-�
0���рJ��g?�W�v��a6�Fs�	��>t[\t������j�A+�VG��)/�q�`|��@Γ��>l�.��3�:7�`�@�ɩ���QF�� ���,J��X�ֵTW^��}<�S�m��l�/��V�"e%�ӽʡ��	<��ZZ^.�������
��K��O��\���`��*�V9嚑c�J�pzy��f�g6^^+ׯ6*j��_MT����*I/WV+\�3�W�
�-U���U,z���рyӗ����/�Gb$?��_v�<�)W�	b�N�&�>X���nGC~=2 Āx���裏׫@ 'Rz���&����l���׿�6m��3g:>�ÁA8�&B:��Ch�R*& ��siK�$�-�䓆G(h@�j����ej�r��R\�4A��_�Ư� TKKT늿
m?�����+'o���yk�j�\�%��xTY�����˖�V�{��.�`VJ�X�a.�f�S��*uM�,躧C�V���8�$r�+��b;	�_�*qG�sy��:*�%�'(Qg)(H{9h)ڋ&�o�p��)k"���9&О��|��,�TF�i��l�}��[y�3���Ҁ�y`���|�D�$�����GLf'���[���SN�S<��u,b?ҭ�wi'�;AJK=��"�MX�iP1Gc�?ّ����	�ą��5���4���*��x���B� f�n�U�'K�i�Z-�k��SE�ӓ1���C���XLE�`�ڥ7-��R��aB���,�1�O61�U
N�4Z��+m\�����@�Z���S#��chU-��
�l�8>�.���s��]�2u��\���G1I�oh?���`�6k��X����Np��_0?֯��5����|�O>��{�A��@�8#�i�(���*��b4r,��*���<ΔgV���Qix����j*>ٟ�)?��L��&��\�^��EPF�|��آ�E��DI.@�2���O�s�i\1��]D�m.4 �:������
-����r3:�%BO^�N���1�h��� �K4Rvƽ�����~���53��X��<������iS%G����f�Z����y��U(ѓ�Bpdꗾ��e9�?z8�xz@��4�k���(���ߏ6�ǀ�x�c�����֬��ЈUn,�� ��KOʖ�p(��d�≅���Yc� �6�aȀ0���ip�ӽ��3u���o��	��X���ɂ=��]�N�@̮�eV��|&C~�^��%�ُ@�hq��;��e�)��OR��b�s��+�rhV�ќc�z%FR���\�T���F����W�Ҁ���^��F~��%z�=}J99�푁��:g�l'����'��/�6��k��X�0�W��h���.�K����L�����{T$ay��1D�T����Z� Uv�#ϼ;$��li�g���K����A����(b��W����a�����
Q��{�E�P{�@;�2�Q�O�,��/	j~��s�ݬ+���5:��d�{���$� d�+�B`�)W� [�)�J��QG�z���b�x�F� ��y�J I{#�i�m($Z�4�FcK}���O��UZf3�P��z�(�d�hB�U��n�|1/���E�t�`%��c.U�	8
����o�����n>;r$��j �P̲EO�]�>����ˠ0�gL�ΡΐQs��`B�m]U''�β�H\�6PiZ.�a����x2BV��U%�(��a�M9p4|O��F	p�&u��6L�m�Qzp�������^
F��y��-Z��4�*�!�MqLLgǂٸ1���9�T.{�[�[������>�H��F'�Q�ٳ&��W�;Gs ���:�~Pp��w�\�ɠ
CI�g�tt��]|�����m�_1<|�=��/�c����jp4��MW۩\%T�:9�L,؊�,��X�(m�FEK�x3?�s~2�����!XV����Q��V~�=��'�r%��t��q�����!�J���A�,���HMhz��x@k��0��+���υ���V����!Пj�������>n�o���c��ِ�����ޥQv�iS�����`���	�9$}V����@��v���sf���f��J��^}2U�01ԚKM�Ϯ]]�S�{�Z�O�t��C�baA#)�d�w"@n��YH�G?L�9!|J��'?i\yM !�:Y~ҫ'X�A'i%h���� L��Y!��}�ר�rz��.]�p��(K~k<��?	t��w><��C:l���'�:�3�Q�����VS�9���J_�+;��ݱ����A��#�	�!�@�5#��9��??����k�&q-M�s�S嚡�_�$܍+fz3<�m���� ���Jr7���7�A-�bN��5�̈́�]򣽼� =��d�FU�l�$���&D���y�H�;ۮJk*�I��fD�I��������O��l�$�@'p��+��I����TVs�v�w���O9��TD�����>5n��o����u �`Z���ԁcX:���sӎ����q��v��&D�l�?��_��I�T�/�=Փ51�5T���b�L#���E��֯0x��ؽ�>�N��P��ф$kC�h1���x��"��'�J3�+!BK'I˅��� B��P���!X��f�����!��	G�Ȳ�f����℻�1��SRV5�4Y�h����l�f
�`"��=��O.�1�MmARz%�˴6���K�:�)T��AE�Q
4?�T~���s��g�#!�� �hv�}��2�����ř��`r��	|>!M��� K{��r\Sc�ȣ�Y�G b�7��\p�9� 7K"x��s� ��;^L?y��|�h������0���~;��l=�>G�XӚZ1u3���0�;HO�i�ȏvL�F&$�/��EbB�ֱJOR�yE^	U�8�#P�l�.EY�������LIc�;|O� |o~ �G�\���~�)�Gh�mKe��,��h����y�Sک�@��={�/��~UD���ׁ)Oz��\�Tw�C\�p�T�q���|JA�g�R ��ŃV�X�:��$Mڗ7�ϛ?�[*���~�+w�s|��	�V�r ���e�2�n��=��W�A��������40B����^p�������'?w�}O�5�g�	�����)6j��W�BMq[<��س�����G
����hcO����R�>���N-�a��J�ex� �g�D�'*U�~uuQT^�����x��H%�t��>�́�M��]x�_���O�����Vn��ǈU1yι���c�VN�Y�)^�����{a�t�#����������Y$�/��O��r4nz%	�%/���� ���(��S�T�Vi��n�2*���G�-^"3C�n��uww�Y��Ƹ	3��ː�*�����f����1��t_rI|��ߌ�'Ĝ�g�3\����ԓO[���G�(��k���0������~�r��t����=�O;��Ҹ�λc����q4�,l�Ǟ[�}#��R�<4���� t��_]J+���*�8*����fe(<Y�!R���#��.j���.^�T'+)A�H�DC��jSC<��"IE������I�_�Q�i�{�~)���q��~����((�@Y���g�{PکDyKTvzkni�v	,��P.�Km���EۊJ�ٯ:����ƦE�E��Ҍ��{��h��V�&��vIT�Z$D�)%�d�<<r�Π8^B�sƔ;~FJ|@V�?��?�1cF{C϶���˯���/[���	�ŉ=�����(��t���⪫�<ж���4�!���ܹ3��q����q%b�����<�˅�H�+|�ů&4�|���OL�S>�BK
*�$�I�S#�Q����g�k�ؑ1~��?a|�?��s��G�52��C����rC��a���T"7,��QG���:]E��ur������`�.�,������ʨ�ĳ��f�e�|�3�Jt�!�X6}Q��D@�KAp-V'��g�|T�h���!�Ż�0+�AWO]�#_3�����*@�S������ȶ�f\�&�<@#x��L?�& ��`\�f��&{���eY_��K.� `�u�Ѓ��v=�c��//~ٶ/QY}%HiCʱ 1R�#\fMv�= Vi���q�=	�����0*;��$��1L�q�O��v7N��#	�a�����w(=����̯h�|,�AK�fx�9A�1ޢ�$d42{��Ҧ
�;��\3s�<⧍X����a:U	be��G�0o$b��fi�6�Hؓy�@���rVuoA�?�������+?�mΟ�V6b��D�(�u����ݻc���)L���d��^h����{� ��׃�T�0�;w��*��Ω�� �g��ء��G������xιN�D,H02� Ȭ�^W�0�˽~,�ʗK5ݶ�9�U��iIJ�p�a�}���V4��bT�0�E���S	,ﷱLN!p::&�_(3CƂ�w�:5z��}�iT��u�Ω�~u�@W�>N=��̀�n�`�uX��MM�tN�<��x���nI�3�|��r��B�T9�r�����xt�⋋<J����lٲ�=��ګ4���N�ea?��;@}0�i�ԩ`^�#��[ĜD��oAO>�	���?W\q�͊��9/�l�K��j\f��T���P�N��^��Wy\g��44,���JN����1�N��=*!��
F�.	h��'J%�LȠ��ahS�%�V Bÿ}ׁ��������#�Duc�&]�h�|:��[�����T��zE�%9տ+^�ra�?��)'^ �hP���	r�v2�J��?BJpJ�S��6����q�{l���s�W�\)M��'����b�r�)�ƌ'����_e�s8\�X� ,�� {`�M��=�δz��7��?�q�رS3ȧ⮟�������H�;��&LR�bb��eF�q�̄G��4J�L=�wͭ5� ��
�rϓ�f����&1U
�I0J��PudE�B�p�Cr�-w(���VY<���i%GUT�$��&���K>tW��������Ph�X�R9D0����S>��zy�9eH)�@'O����S�V�%��@�{����\��.B?���+V���lv)͒���ʷW��c�?�D<��Bc�{�5��>F�9P�|X*Ü�e�}˓�'�H�0�W�px�y:s�����ҥ~E���EXq@�^]��f�8@;�p>W�89��U��C ̢��6P�,ib�n�JKzy��@ί�;1L�W.kl?�R��x݈81�C��5kF�[ZQ���L�D~�DJ�&7dL&
����yɈb�NK69���ٰN9hX	*�s��E��	�*�
���(�6P**���M;׃��(8]sӝ�:�:f�tM<T�rݱO#������H�����-u\<�Գ~ys�����た?�x���#�H�_�l���Cp�s�F�����|�l���{ M沰w
 ;V^n��x4;��b��a�'v"\��{������}
t�R1"���n	")7yǎ7}�C1x��ۆ�*�!���tV���b��229�Ә�^��bvYaz���Ri�6	�?{%��?ƙ�{����(.%el5�XI�0�C:z49T�(,���^��]],A�ͫ�����݅��,�)�O��z��T�?����o��4��)H�� ΀y ozR'��oKC��<��Qi��+rs�\;���Κ\~�bM�������H���e2͛ �q$�m,R��=���%	R�.��9h� F�xw߯��y��y���������?�G�{9[�Q43�kܤ��ɮD� ^�(�m'��t)>i"�[b��+O�qr�d��������gz�/�P�;4!Le?B1���}���0	�/�xc�jƇ��KX��v��]��~�K1{ZW��>Q���U6)
5�(V �g��6fդTvH�>5A�*��*��̴r�Aiz,�B=�:��Oě��J��S�u��+�'T�6p>�g]�'�[����������4ো��Q��Ӧ�_��?*4�<,$���I`J�f'��� l^��f>H�ll��<���K�9�?������?��/�~�F�}8�tr�_�H�G���e���ֈ��T�6�g!Jo��4n/�r��ꊒ��Wę��-P<3�NiђR�����Kq�hiɁ4%8
�\r�َ=��R������0���k����3't�G���"j&X���ם8��fK`2� �w�x���2�|��
����M�x[��T�BZ%����/����Pcv�D��ai�t�|��.&�)#BK�zG/]:��$� U� ��;��gL��|�K)B�%9<(�����r�0�;,�w\@RP��Pu��x髯�W��u/���a������/ƾ��h���T�L���y(�{j�|�G�03q �����t��Q�k2�T"�^4'.���Wx�� !l��e�JIӿ�ƆX���ݶ�B��c]�U9C�o�0l٦���w�ʨ(팡c�GOI��aq�%��Ff�@�x�D�:�*։�~U!�ȤϻҤ���fYO�}G��^p
���Р�Z� �pJ+^�J�{�eFHaX����6�	��'�9��.{W/�#�bn��U5򶷷EE9<T?��P�L��� $^p�;v��+�H��|��>����O/��� bB���-��m��c��	��b6gl�v-Tq�9�n%�4'܁�~�4���c.����g�5-���G���NqL�T�Z�]4��PRTK�����E��P	04�=���A!�Cf�)���oեp(��L��~�H
���P��C��*����pg0_�R?.�ւ素�}���țʃ&9���-�2�q�-H�hDS9�D�s��<t�������%S�^������٬y+����+
���e����
'����K�ʾ���t쑄�/�����������q�78��k��=����������0�پ�2�����0��� �����H�e����J�ܮ�b��-z:Kgd7r��I1dH]��7@�%�,���f~'?��qI�����Sy�N��Si����S�:�㭓�eiq��C�]���y]]u�N��{���'E���?��ӯ���=?���G	ay���D��`��Ѯ\\p~\�uҮe1n�x�$���^M�;on�}�91��	��u�cR��H�^>���w������?�{n\y���w�;����΋Є��=����ߏ}�C�O}*�.s������U�A;�f'���N�W~�R�S�qS����sQl[�{��سm��|�3�9
5�C���*��6Xy4�N+;
"���P�%;�����A$Y��LA�n̛,� ~�]��ɴ�Sr�?B��DxR<�SWH����s��,�M�nE�dL�C4�"w\�Gq|Op޼yq��sb���T^����ԙ3���*�^���?�C� �%��-���w^�u�]�| ~��~ϯxL�4)����{8�jٲe��}/.����4�A �0�k�&����Ƒ����bc�Ȍ� II$H�F�����O*I͑56����;d�P�ɕ�K�J�P�)��p��
��L$͚��wT�E��%G�h�L<Dsr]���I�^h�?g
��p�ꕼ�~�d��6+����ſP?����JE�pYIEz�-)i⩐�s/��֤�S������(g@�ɶ�3gN40;��_�&A�3x��j�*�?�er��f������+������ �Q�y�>��Ұ���/�&	�fw�X���9qf��-����"����+�v;�>	� �ZIˣb\�j�e���(P�7r5��%�-�YqiQ����P�6f������R�I=䡯r2;�}���Nq)��DY��ɰ�ݓ  K�{��[6�d^ѕ/�#$$Ɲ������+�
���0.�P�"���� ~�?L��yR��J�<p�4�M�6�_�x��Aލ�����7W��U��,G�'v�ٵg������p$�����7�����}�d�*�1
���P�W�-��l��#,� �9>KkPE�+I�3�<����6���0�d��yǖm���
��Ͷ�]U�rp6��uy�Wג!	��Fz4fҖ"-��k�R4�5��΃�O�ד�O�N��s&O�He��N^���t��nܙS����J�#t�Ic��8�#+`R�ڑG���c (���ϫW��A����@�''*�+<�{'���Ė9���=n��6��2|x�Vnggg<��36�pr������o8�/E#X�1l��U~���&�˽�?~�,V�@�X9s� �;�:���J���qS4��+<�I@$X�gwQW�68�_Ti��O�p)$�Ř�<L	���a��}�k����	b�<^�>��r�����ܲ���]��3�y�yάʚG�b|�Э�� 4�-*OĶ�!���Mc�<�[iDE�@
�����9��y�;�������s3��J��y����w�;bŊ�+��bE�ر���"�[�ƪ��0{�SQ�gyȗ|tX+#sRg4�C�����=�o����|��^�`�])16m������{��ų��,+;��ʩLi�e0 ���}��}x:ǀ��{��-�\���SA��]��&m�,
y�UW�n����';/�� ��2��P.�OgW��K?�Md��SaY�,�I9 @�A��l��v<��VW,�Y����`5��W肁\���~�,XJ��'c��<���s�� jN�5�΄���Qe�T�D��)�.S>��/Y��p��ɲH佷Ez	M�;���%�٭�~׮]�R����fg�o�:t��ٸi�1��C�|3���Ҩ�������o̀|��fGB����K�����]w���3�|w�y�p�v��7ǯ��:]/���yϼ2v>q �j��_����I��������Y�c�x.U n).	�z�|X�O�'�َ����9��C���rLsQm�[;�\�?r<�x8��4͈�aLt��x�Z갣��f���5epq�2p�g�z��RXly��_q֪8�H����Oi�7 L33�&z��м�Hg�揥�,�Oю09�l�(�^o��ظve�Fl6=��2:f��b���^�.:�k��<q��`X͈�|�����T��^r�ŧd�LO��-[�������o��F�y{*��*"I>��$خwS��z��fNs��e�9ȾO��[n՛q͕��O����/X�Mٰ49�%[�k����#ќ�K��W�*Q�/��W
��[��9��#�ϥ� {@�6[dhB��{#x��IۢQM�ڋ�l�$�K���D���%ԓ=ɔLx�H?Yz�UY��._F�_�UH��>�2>���8��GxF�[�d�v��Fv̟�Ȟ�S*����3;�I�R�����X��_���i-o����O^�.���߽�' @��/�.S���p5*�P�:S*�	S7N%����|([������S=и�O�M�l2U�8��l�E����7?�s�n�U��͇�~;���R�-i��?��������C� _��Z㡳y Ԍ�l�|� ���ʯW.�؛23���t�萊�R�܄nѥ��z8��gz�O�mfP�^��f����+�썶جe�C�1!g�F>��u�#��]�=^�oL�}GA�^P��_���h��ʞ�·�P�w�s�s���:j-S�X#|������7��Ei���z L�TY��t3�9"D�-Z�}+X�����D��<�L��z����P��k5:e�c�6�����(����[1}xw�[���(9���Kۜ2���7�j�����Jy�����X8�*ХPY�/�ƣk��J�_ʬ��&�W��։յ�[�O�L��#>����5=�UW9)��}���TR9����{��G�ˌ��w��L(����>����_?�T�,���DItX��5un̘�j9Uh�4�����,RI�Ϝ�i�Zv�U�u�����_��v����|��h���
�A��h`ؘ���	��>5���<�g�~�u��G�(��yꀌ� 5M2d�$wE�3e \�Ρ*��t+N�
��g�� �7k�Xh�/APg9��eJ��|���W\������g�Q �<��t ��C�K�$���3������_��V����2���W\����\1�N60�y贓�����t�"��)T���+O\S:3��K��<����$x��`���M���u�k`f6`�#��_p�5�E�7R�ٚ�{օ��l-��1��r��;�9�G��@ȣq�I�	�}?6!楁�u0�
��ҩW� ���g_�=�m� E|�Q��4��4�ʑ����Qf=���&�O�����W^y
�0���}i����&�N�_� �o�Y4�L�T�%�����[Z�
�i`��K �z	��'g��t�\-RӪ�i��8ۖ+�z�kX�0��B�c���\�B�Q.�G
o��1!�_u����t�}|ė,�k��Қ���y\��!r= '[Ԅ.����k���P���$E�[F��=ݬ�YB��_1"6����cG&�5W��}��,�̎u,9`v��֧s<[���={������c��S ����&ߎ�����︷���	a^��*�.!�q�"����5�B+�x���f���ѵ*E� �)��p�@�="�Y�i�`�Q ��������_���|u&�4!���l�/ ��C{�^ @%�A�n<�� 5�f-� ��4��|�?"��#���T���p"�H<{ �#Z=�Aϵ��-�;���U���'�']��|�eۤ|�fڧs,-��_�奮�%�_�}�q�~>��w��
�o�������#�|��o�O}�S��vk׭��ߘH�?�se˱0��k���~�����^6��)c^�����mo����ߍn���~^��8���tg�K5`���gg(}�~LHi���G���iI�JӁI�4s��9����ӳ���J�U�*����є���������	�R�[�[�&�^q��`�^y�MWR.���]m "9o�"?�Ϻ�����?=�Zz !?�8-�s_�SƟ�IZb5�,z�P�% �.ctǪ�W��Q*�R�֭[�z������x���h���E�U@9����O��۶�;&��6�'������On��6����%�\����)ɄH8���%�[#  �Z�C����%�	 *�JI� I��%����}��H7ދ �S�R.�!/��n�4�%2����,��e����4&���5e�I/�Ɓ���yəN)uaZ~�����M8��u~�,�䈣\�#�2�q�1)Ҡ��"e�\f����Έx������^�2ۿ���g�MQ|��)0����F�0f���/ۄ8����d��p��g�% �^aO�^��Wy�_��_�w���{��{N����
cZۣ�>j`ONNz��S�$4��
	�$�$'8+?���5KD���h�@<-��:���Efl� ?q�%��iy����E"K|R�S�	��O����^ �W~T���u�/��,���4b�+SzB^:9��)=iu8�g�D]���@�W��<:�?��L��u��:�9������?�q��%/y�����u5,�����ـ�0X������<��gr��`@ǒ�3��+W�w�}�����6�h_�q�9:ޭc���r���!� d	�W:��3�%�4{@�$Z��=���Sp�I�I6�*�g�
k&���*�y�}�E~��^����#�#<�'����m�$R�	^�.=g��cv�/�b
�`2X[B`b�ͨ�P�Ӣ��-F�3���7K�
��e	`
�c�̫_�j�̸/~���
Y�f������ �gr��6���S�����O�x����s�E!Y���N��{g��=��uu4�e�Z��`,"��*�'�Sb��Dc�~z�V�"|Pd�R�@@��!),s�*��-��`p���T& � {  �^��0�Y#!=�'[*��|�;O�8���Һl����>� o�"�z�#N!nМ}�3xs�O��Fg�܈�8�L��4�/h�#t$:�c3?zaL�w��65Y� h9� @�{Sk�f��Ǵ@+�u�]��vOz#�]��GӻmO箻�:�������{/sZ�'>�	�:
�iY�X����~6��d���V�:	�/�/�ϗ��M�XC�\��P�ܕ��K�HҪ�"̐4�9@A���z�c�6��eV ����gĽ|p=�gq��po�K�Nv�y�gh���(�����L�_&y���!Oy{�[���}�o�8,��\���T�'i��9�w�^�ͮ��jۺ�l#��G�W��s� ��8��1S����>'VO͟p���y5�صO��K��v�3E��R�4l�~���g=�s},�\�v�[�G>�S�&��g\��dۃ��dҶ� P廂9�����6I��Kq�,�7;��H��Tl
����L��v�9�4�l�v#~�z4�c�'�2[���{c9���hi�����#d_�H��_?r��0�Q.ۼĝ&��h�k~D
I�$x͋�x{+v�Q�g1��hEM��FkV��.�f9����N�D �L��U�Y�ȋ�����5�G�q����d��\G�<�].��)5f��9W�2�Nl^2��"4�xX�l�.� y���u�������/u6Z��D���#/_!?V�:3\�.�r2�,a~���wz�ٕ�g΀�K�Y��<��7�é_�/W,1���A�p�6�X=F��v�9;/͸ա��ˌ��Y�gŽPF�J-#!4�1��7H�H����G���)7Sf�Ń� 1)D���̄�ʑ����]_����ʕx��k��1�AD��ϸdS�p��h�܏�����?;`v]߸i����p�����yj٣�;�Xʧ�N��K¶�%�B��d��Z�*6Q� �Ӓt�齰���{� K�^)ܛ3���x�n�13���oz������ <Z��b���s��yɄ �1����%*7gz|�!p*�;�UxJF��Ӳ�M��izxd<1y��D_�Es���w8�<��8yٻ����3W]�1.|�����Ȏ�ٵNK&�ߠ����i�r����� �o�ѱbl,^��?�os?i-�>�	����~da�)7�87�����=4;3�q�+�7L��0��W��e��@�~�D�0��7�!�B�h*�H�^��AF�F�V��r%�����ԃɸFG2�2?���.�����Z����#��|�C��V�NԼua> ��8��tF �ㅖ��p"�=.���=qf^�r�&}�[�G�G��� ܨ�cQ�`��R�',%G�ʋ6�����8�=�^�����ݓ ��2����k����]�:����b��+UL�Wg�W k!*pz蚈��I��&�V �	��Q)O�W�*���nVZR���Vf~�T�3M)��$-����Q�F_���_��yY�K�MI��u(��T!Hj�֜dk~�1������F�<>��@��:m�8hdB4ma�l��G�NA��-�� �9��m�"v�շt������ħ3:��/��P�����l��?D^]��B�������q��wH�dg�)u�`�g��q��"ux�&dQ��r Jރ"�D�W�a��ʼ��R�RAN��@za�nSA�����*4�@'�/]+��6�ܱ	�G�O�;��y����R<�S](��a�w�dԦ��k����Q�K9��#�%EG~ܯ�ۍ�?9���Z'��2Ҧ��&fI)Z�ꋷ������8��L\6���!O�i4Nf"ѽ˶f{���:�.��c�1�y�) ��7�??����u���}J�2��7'x��<��)��a?����k
��rE��M�4������J���� �<c��]�'O�Y������`��T, Ng��@���_A}nNv�<X�|�J�@J�uq3�\3�A���ɋ��kP*H�������7P]�,�����?�g��I�yz�$=�Rμ�D���5�Z&�5�3�oǽ��]�B:G }bO�#�E�K"����@Y��WF|���ěR5��&ڟ��) �}˛7I�񙨧K.�۷F<��Z=���d�.�h0⶯K4���=#��Dn����vo��?}�Ψ�� ��%�W��UR*O< f�T�5�j2�D��S�<nښD��M���kǉ:+�E:�� k�>�"�p,,�Sr�� M��b�щ��D_��6����P�;���iB�d/4�/�=9�`R>�E�4`���XU^˄F�8�
��hđ�O��i�Sp��SV�Ƚ�� �G�� k�=�ʣ�Da����tՅ���vf1gr��^xI��ֻ|/��݇6�E��,��`,^���{���xͫ��G�/���I�~JG�j����F�Sy���2��!z����{2r����{�5�E~�"��]��{c�%�R�&r���X��?��_�я;�S�_y���=�F�Aaet�=���I�Z�8�]ʋ�B ��&��@�@�����8�W|�-��/-�a����}�_,x}M��O���P�&���/���Z ���S����������8���?6]�"��� ��)�\���� `>1З_PY�� SEP�͆��=�@�}�����ň��u"��g�\g��Oiд��Lz��i�\>S�(���F׮˄�s�����9e�0s�6t�����we!gr'�����pt�/��=� ̇�=����b��c���F��E��/D����qC	eG��?���_�} '���ky�_��ȭ^�?�p�~������E�@ ~���⏽>rw�0���7�R�vz������`
�@	eg����2���%`n"�W���g��>t�,/���5���p�VcC�a_i>��vBX��� v���E���n$ppr��xho3��?�A,�>~��۾��Q;>y�cH+�s`vZ*�2�ÈQ"H\i4�?m-[��Ŗ���Gm�[�ŵ���|T��S7:K�F�bE���=p��40���2��?s�5�y|a��hwә4$w"�~4r����v{t�/��#q��q����G�k��d"�?�#�;��+��x*G�)g�?���t���gp)�H��~"r�_��ϋع;���l�g=#B6t����W�gp�aۗ�W09U�H�=�J�P�6��V���D��TC��w��W����"�
ȗ��T�b�$� �r:��_hX�t�C �#\��=�Z��:�o�K��2ڔ����(%�q7$��B�W�Ӏ���tZ6����P��ß�R<��7�@>A��b�b���?!�L��g��5X��f��y������е�obd��x@�����o�I�F�֯EW&g�/�ܿ��p���q��ȽZ�o���&ƱC�]"�3:��������[p��Qt��А��*�+͎G엽����>��S����Фi�F�Y�=�%��\%�4ed1�H��z��T ���y�-��$V�X Kz�q\`�0�V�@XZx�T�[��Q�4 �ɏ0���"��bG�K��0z���S����8��I�
h ����x M��0xk���!�n,�����"]���:J��-5v`a��2�hT�S<��+F�$���ۥe�F�Dnպ����No�Y�D|F�9���,��q.��얏3��;GdX��\f����z��"04�m�G���"�̫#�fut�z�u��u�tsd`��.��S�b	&@N.��&�R5�,����X)�o%M�_i5�j��Yz�&���>i�4�4"s�t�֖(_�Lߝ3���^A����  `��[P>���m���뀊/��Q �����l�Y"b���{���d�c����+�u�uE��T�\���De��H���"N���DC>�3��աA���k�9i�h��+SU�.���ޑ��s3+q�ʧ�T=�>ݑʑ;}5ڦ������VqP*�7;�~tOD�C�W�L�H��ء���5h��08r�cQ�Dgr�)P�R��I��*ɥK*L��J�ӥqJ����sN4���lF�B��E���z6�8.2^F,~+[t�*�,�,��/��b�Ɍ@���\*��{��g���
l��.Z��PH�m��J��  ˖�lh�㊢��=���E��Ӡp�V8'����K��(ܽT�8���d���"�4|F錇\�Fn���{���\��#2�G�+_�_�!u�����7"?z�EK5'�@!�����\ir�"W�(�]���to7����c���O�:�g-������U� �ת���Q���Uq" �wi?�YZ��?%�C�\��~�gQZ�,��I)C���2����a��6"�k����s-����5* inضѶjN��ܲL�hg��p +�Q~4��.%�dR),Ӗ.��+�N>��;M���ܞ�极���g����!3R�9�-��)�7\q�-���G#��oGW&���?�����~����xjOu�5�j�
MP��d'��I��ֻc�U?�׽&�o>�Z�t\�������D�<�Cv�
m����?κ@ME��R�˛lhQ:�C�x@�#E:,�Ti�;.(o�I��	�m\ٺ2qdA�
iJ*�i��F�.Ҙ�#7�b�ظ��Y)؅J ԁ�����c� t��p�S��R� v���&�b?�,J�:��O�2$:����=���fgE�a�t����E�mgW�?ñA��;#��">����{i���)�ǡ����0�J��)y<��N����[��K�LIN{�,��_���|鳩�O���8��sO������?���ۢ!	��&��1`�EuR�T�~ĔI}恩"���2�z�H%Ҙ�K���� ���/{��E?�:��N*Bw��⣇��������*_���i.������D��qTm_'�8ъ?��?��{?o~�O�e����?Y�ِ��� �-)�A3���m	l�7��t ] H�>�DB�ɬ�?O����?s���۔�Μ�v@bt�4&�OjN��F]�4(8$��ǅ��().:��������d䮖���8W�����w̑/l�]֙,X.�jE��h=�r��Oį������DC���9��0vo�%WH>�7;�VbS����L������	�괦^����yΕ�ʟ���V�|i��J<�rљy����f�4,��	��ż�&e�����9ى?����������O��?�����7�q���tp�t��߯��� هM�� ,B�:*���7f��0����G��~�Cљ�)8߹~ܳ��u���L�KDG���gp�k�P~�_��Lp��+�#��.����5��=	�g���N�����ǯ�u8��`j�n�JE^0�$@�n�Z�\Av`�klH��>�4��ǂ�V�%��R4��k'�uozCLl�T�5E. K��<hb�F4��Ё�hN�T�#L�<gC�����,
��v,�[����_�ۮ�.fv��|�c���W�j|�����ۢ��*pʿ���M��d��d�Bt�z�\����r.��>��V��#>ӢН���d�0�oq 	$����;-5
�DI<7*9��`�$)�$�>������~(֬��l��2x:>�;�1>wíѐ��N۝һ�Xk$qc_Z�r�G��� l�ELc�-�-�mT�� �G87j �3V-�������d�5��#�hb��dJ̊��}�˱���T���?f��:�Ri�P�ks[#�咴d՚�RQ?�Dj��(����1��K�t"�P��M��Y��,pf)"�l�0�Do��@�f��Ā�,���) ��D��}�W^" 胱f���O��\���&i<*��Ű�\mv���p�pd��S`�qΎ,��Iy)��)*##�	�G�x�[(�c����I/�P�?�F���8���X���b�uR�TD{Jc�Y)�Y�����&_d�y�� ��<7k|�Ovr?~��Y#���9c�}��wQ���ՠ��"�|(���d��_T<ZREU�*� oqr��}�g���Eq A �s�!���8�$�'����5��e0�ζK�K%)��eI&"�BNV
�S��k-��[��,bd"�j�4ٳkw��!Elp&���#� 126�rU@A+C���0O�=d9+�Y�İV�9�E��}���A�����y�v�QãWdɬRvb�%���jӅ#"��wH~Ī�2�5�Y�r��C��4�SX�Oe��p���-�-DU�+�B��3y�dϑ�_.Ef2�aa�Б��y-M�g.-� e:3�q��������H�Bc&  ��a������DC��2��;O�rj����]��R�
4�^�z����v�*����q�Y���#�f$��M.����/!���̇�ȳȥ�(>)h�F��Xv�, ���{�}a����U�	ܒ�EtJH	�@�����y�`j�9>��tf#����X�����T=rH�@13� �<� �J*plx(�C�	0��Y�Y�dl���Y�]�uS�0`$��r(�Tiv%K����V-��y:h1K��4��sp��������h�xRhy��<�����!K�/�'WLƏ��uEwT�K}��{������I#�$L*�R�4�+��uF�
���i���0�`^3��.�&���/��L#��~�ɇ�-#8��إL�.vQ���C�+y�7����{� �t�s�� DΡ�AK� {\`����L/x0�fZ�a�N��@g��8�c:��q�L�4���z�@�pq����^�kV�ߺB�����2XNB��1��OV��ݵ�e�8)�� ��x�ZBtvu,%I�6�^�F� ��f;N:y�<���72_�]X�R�?V�Y����.8����t�<k픣�R m�Q�I�{e��� 0�[�]�3s�s��TY.k�z²�ih�J�b��TEC����#� �����g�˙�t�[ ���(�6-��;�9ZBK���3+pX�� w�dˁ|�����<�:�Su�������E�1�J$ `������lT���j�*��ԍg��Tw;�����,:
%O�*�Ӳ{�˞���gt=r9��&	����I':�7��'Ŕ8������S�{�\�8gJ9I.�K{g��B2�s�%Ĝu���k��P$Ta�U!TP�K��4�����.�IЦ��u �
�i2�f�4ؑ�w����;F[9��2[P���idt$J|/Y	!K�	`R���P�3'>˃r���s>\ir.q�/�O���@��o����nyqؼIPL���W�Wf�����y�F� ߃�$���W&��s�`�!!	(Ś�[�
'a�&�t�~LZ9%�zK���*� h��џ1�_���ʩ���ck,������xd�g�cd|(��V��"ś<D��W�t�E�����˛��`�G�u�M`#�����Sn��rO�w��^����e!�W�7��Cg~��,��a�3��D�v=�0�9z�>G��΂Ah��'��
���" �Y����P��zzBNP���Sٰ�WF~t�i����FM�G٥r���<m���,&�+���b*�eD��Y(?5��Hk�G���]r�h\��+@d�)-�8��Ίa�,M�ݷ�������ipN��S��+rB�*����$_��]���Y�`�)�s�-}+�l�N�w�~K<��.��k'I~09s�?	��X��/�o�2s�[��QI���+!�t�����y�*F����ػ琎��g������������b�c������I��s�i��������y���&{���
��X���ĿԬD%@�v��V1:�h��ڸ�i&�&K�N#���u�+-.�thn%�9ж,�<��;��[J����͞��/�0Je��X^�,k!���'�����/|Y�?��f���VU_v�d|��B�*��ȗ��ﷂEG�j��K�Q��gV���%C%i�BZ�C+�
��T�����C��Z&��%�9;O�_瑅a>�-�t鯊VˢS��I�.���`!��\'3��s�C�0O�%��,�Q9�s&�wz4c��^?�J�g
&&��:-ɾ�l��r�[R ��('�����o����k6��3 g�e"9�.՗/�1!*ד��$���\�M��+�2��	�*��4�:�g�$^��ϟ����h׎G����X�O�bsڋs\<j�r��߀��9�AFʛ�1Gls�^,�����>�V$^���)IVfV)7E� 'ރS���j��C9l껫Wz������_zȭD����A���G��sؒ7�^�9�|kg�q��n/�V�%k.�x^4�Cd?���8'	"�K!�,tO�f͛�R��V5�����b��T�8[�REֶY�d����s��4|*�|:{�l��oV�%���'-� ?��Hᒍ����R��Z�L�>ŋr;T�;邒�'�.�t�<2'�����Xڝ*O����p�`9W絝L�,V ��~�+ �:���hH�gM�K���2���� �K$0@t�$W:�y��j�V�G/�e�aP���X��tt:К�	~���ؔ��4�#���K��2A+�R��hJ4P)���7�9P�E��c ���L���[��-�@pI�/�[��t�q��t�b0;	�o'R9��"Iݬu,�.�Bw��	����Q�����(�1|�J|��k�{�
`�9ޢ`3��7��G��P�6�鯝?���<y�^�J�vUn�����#`jx'!��+A
O�Ư�:�G���C���p�'�T�9و���y{2�Ѹ��?��w�m%���u�^���$+�'���\pH�9>+{r���-�Z'��vK
w���G��bR����I�Jt҄hDW���\)��e�T���t����?���h::�;NSa�A���(����t&>���8�-�ގvKgf �^H3Ww�-ž�h
4�[���f4��h�^oD�V�_��ķג���|3��9��Dۨ뺮����oՉ��S��5XS���j�v����̐1��d��j6U�� o��wVg!>����Љ��6>_����DM �����Pq���8�H��[l�a�RN�(j	�ֻd�K�O��9�)����3��|)5�Ӛ:�\G8�~�NNe �T�JE<y�1��Z��,8�Q?����M8� �7��D�2H��0���J��|D�Ѩ�)*��g��i4�Q:�Ĩ�GC�M��3.?/>��������Xh�Fna.��RT<-�\|��wA8!�R�0��45R_�9� ;nq��s+�3�����]�x�s�~e��y�q�ȇle�]iaE�i4h��}&Ne�$�\:<�C�L�I�1�#]�8�qj���_ѥ��St��(JM��H|��@�]����4ě�6��t��\^�-s��ס8'U'�:��{Թ.�ߝU c���ctb"�F�ew�F5c6��x�)IOq����bI�*9��nI�)m���+C^ϕ���P`3ɠ�/c�!:�h�(��&g@q��
�L_����Y$�(D),�M�ud�C���I�0!,5�c~Yᾖ�5�)�������
L^�N�����Z0Nae�9�F��&:�Y�5��X�}�Q�[<�M�H����d�9�4x�4n���邴Tq:vߙ����,�3>Q�a���E�[�Xg)���HG$���%'>��ͪ=+R��`
���?him� 2��l��ck����0H�4uv��~zg<�'��eQ�)����{�@���b������\����/0Qq�ܘc��*�X(��$�U3�~'LvZ�������`	�ƁR6X3� (��h�:W�U�(8������X�d�:2��9��"k2�!E'�t��+��ѨSi�\�TF�1p%#�nк�P���d��=>���We7'���ҥ#�y+73O�P.���R��9��CK�
˔J���p��Ysؤ�=�X)�w��,qVWE��Z�
J�u��u&]�_��(��Q]�x��/��� �O�?ֿ��ƼMI3�-��a=\��tO���art�j}�0O�ɣb�6��W.�{aL�eSn�y)��4�K�%f�/Kkzx:,M	��<uX)��˦�<��0�de����hx���wgu��l��i�Uϸ2>���]�嘫��!6mF����ѕ<i��V�k4�4���l�|;4�tME�J	����ƹ�,]�Z$$��I�Ov�&_b��\��e��M
2��K�8�u.�IQ��u���ֱ�g��?��O�CX�^��)z�C�: �;�2��S̄�H��:�N���@|������ش�B�/�K�;K��,^�/^��6w���s�(ТѴEBtŹX�`%8k%k�bv,�9�"�)(m�0�M��_aY8a��G�q��D�|�>��!gk&i�_Ω��ɎD�҈�g���5ͩr�r���tϦ���� �wYIC��^YЄ�{�4y_������/��С3ߘ����s1��tW(��{P$���2S��{Ё�����,��f���/��O�����p���x�$x*+�NV��=�Ԟ&��4� -˃kdj�4}�"�a�C���`.�h$k�L���G� �p�I�j\ �A�0���잦N�����GJ1Ht�0��AfS�`��B�$*�!�py�Rà�"/BS9H��%����} ~ɯ�8)�$ �!K��d�����������_��_��~���}ݲ xn�D���^w=z$�Fǣ:@�nd62}�Z��V�+����#K��_�Įp��NO���p�(>��^�h1*�}�<��3F��	��z G�h )nT�+��Դ��݇����p(
ZмhM���_��@-a�d�e ��hSH<U6�श�Ad�n}�0�@��%��?d
�4ә<Ċ��+�������c�N7=�q?��F61R�����%W9n9ݲ �67o�������	�tP�X�6d�VUh����OD�{ƾ�`BB���Z`Ʌ��hs��t`�6տ  ��+�x @z�� 
&�Ъ	D"ro@à�}P��Ԅh�Lb�bvv ����Df��td� ���G�U�o��KZ�F����LC ���������sr`ͯx t�n<�D�܃d�2���%� (�ù��������jl��R�/�[ 7j���~�uq�7F�:*�����w-�vC�HJ~I޶�9l>w�Ԍ*��y:�k�bZ�" ;�:<�*F~�U��u���44oT�H�zJw��b=P���i �`~um~J
/!�iz`��(�ѕ�UZ��k��3/~�U�!̓�K2�/Q˯{�/�$C �p��p:��j���Ņ��$@+��_u�|�}��{�ֵ���|{l�v��XN�, n5��]�����mOD_u\`�Εܵ�$讄	�-��# ��_z��&@IW��fh���M
��ĩrSu��<D˛R��ﶠ L � �J�P�`*5k!�1�F9x܌�<t��S�G����e�M�E���G~<�?�7ǘkj����t�'��H�`��R����z�F�e�y�Ȍ�PZ��� � V`-�.<hSz �Ѷ�����Wc��\��t��N��󮟋O_wO�*+b!WU�U����ڼ䨢Qg�#��k2�Qq�����i��P����nW�<E��hٴ�T���0U�bЯ��C��=��O�hA5�Pg;V�6H�Xh�^����2�R@@C�o�^<�lŵ�t%�� �Ż��i�4��JK
Z������1��G�E�G�
�J1l_߳C���X��˙���'2W�׍(-��Z�n��Ӹ$��X{_�a$~�=��OL�с���TC���> A±`K�8��ȗFtV������J��OM�̧^]>h��"DR/NF��6Z��hu����8����-E3���U���j�Z�1��������TxG�vE���n�C=m��e���&�,Ⱥ�k��T�"���H[-�������s�N�/Z�m�-Dk�O����::�2���!�Z;��
�W�&~��s3y�ي���Қ�V#�j�(��0>�[X�,ʌ�����Uк�VK�Q�@�Mo>��vA�u9Wz��̈�xC�j�|��Bf-`��� X�P�ӭ�C4蒐Zs�[��Ph ��J���s���Ҩ��~�],G'?|z3��_i�(Y{R����(t�.��=��Ovv/o��/(~�����t畲�vE[RxQ���s�׹��RaA`i����Y��uݐ�_�J�e⺭���T�zT�um_wV�W���(�ף�oG������5Z���@7�ʿ%���Љ"<�[�AeP�T����ry�� ��=���Ǡx:�(�_)3�[��$@��2�7�J���X���|<=[�/3�Nǻ1�� ����{:c�� �����?����K�+�E=��<�Cw-!��%
��$+�0������%��<)��$�i��4E.F&6	�ei�Y�n��\����4�4|���N��9I3H�B�0U��):��͊�,\~�'4J�ƞ!��o"i��薭��W�B�+ϗ��,���^�!/������Q:�Q������2�g?[Ūŷdw���YS-Z��-��Q��-��2Q��+���+tK\i~������kV�o���c���7!����_���ǯF�:�.��K�J��~_qH �(N�����`�8%��6�9���3����G��\Wq�A�Y쓽L�D�fU�׵* zK���3P�߈���Q������{���@o���o+'���Lkq$`�����ٷ�|h"-fW?[ �M�ԣ$͉I�ym�S��C��O�d�m/�9��Q�95�&�2�z�`Μ9y��䭟���O��n'ղ�ep[������o�;*C�\m���)J�O�
C�p\�ʳ�U1 ��`�2=����D< ϟ�HJ�pWRu��Ŧ+�,����@�Ik}'�7 Q��t�2�����4��9�/>���O�Li��]7CB�Ф�a�1�K��']Do�?�HD9��a�s?������B�m���C��tR���7 8�x�r*�^͏�}��شz<�����
��l�_�埋��x$�#+�éX�7"�߂K�8*ME��K�L��hD�(���H�[�"i	�c�P��SQ�XQ�y�JG?������"kp�5q�7�(�D���< <���ƁK�sQ&��	8:��)u�$�to��r��׉�IS_�E�`��X����d.�|ȑ?�C���@��V*cl`�A�����/mUoD��������L)�12<+��K���X�q�i����{V|_5�  &	IDAT���)3	���J�`�5�+W�Q�D��� ��c^��4 ��k�i�SӠ��b.���h+��EJ�U�*0=�O��v$��ב�Ce�F  X25zC@�F�x@�F#?�n�]��|m'ij�[��;\�U�¬�����t�F��k�r�%x�ĉ?&QǃX�G*fj@�GC򨽫Y�d#P���V�ܲ�\.J��%[�Tu.ǀ�|@�o�aV1e�(��O�-��T~���8�g�^�Z꾾B*C��b�`n�M�evˢ�����/o����?呵��B4UG����$0c ,��mP��0)Rw��I��	�����.���d�����h,��%�Hz�� �h^@�"�09��u)N�2 ��iR�Ȁ�Y1t�������[�%�k�[bf�J�=s�p4 ���m��p٧*Wz���Ԡ���NS�l\(�[�����Qo�FbS�W|*9��1���|K_I*II���/.�8o�����et���\�wßš���|'�&��[#Hˀ4W*�RM�Ŗ4���x��\8�-�!nL4��pŕ�*�jT�*M�������+�!�V"�\E�1��ie0�S�
�v��@�/�+Џ�!�D@STr��6s ��L<����e�4F�a*���l��@���%z
�=�Kz�Tp�A�9����TΊҍ������T����X3Љ�7D��Y�K��&�����J^�[�2^�Co���)�2�ep�Q�����]a:Mw�u���
3I]�/]�C{⁯�w}���::�Qt�-m� C�Ap $�&}����b�U�kX����Q��C��X�8d�@��q�.�h}��O� �ad��=�%?� ��W7��^w��21��~.U(�����|:����Ŕ\�d��T�b?�&{>pg�Լ)� _0�~d_�6��qՕ�ź��F�XMech�����	�V�:.�����k7\�����n�f!�����û�G��6��TE�my	�֬��L=N��e`��4h�`�5{0�G������茀 ���1�4!�:�k��e3�͊��<t"�� 'I���fPg�gP&`�6g��������E��Ӗ�����-0x�L �'P���f�Z��=��X����@����i۾P46>`���a~��.� �\���m�n�"hf�+׮���Ւ�����}��%����R���-W���L����HlX5/x�3�L�2�e0�?��=�7��6�,����n)���Ե������+�!�i' ��d)ߌ��#~�4]W�(ac����J=�<J��q��P]��wX ��l����8�w�4�Wx��|.�1рt��~5d�8=!48�7���Ouؒ������dK�s<�¯Zc�̆rIZ^�?�LJ2%�j����7/����Þ�Ƅb�4oR�O�R������W��������|-�椝y��|��R���IZ�'����*�_t]as�],����@��ω��_Z����-	�����ʮ���t�2�) J����V$@F���A�%>��Z��٦��(�S����.scx�% ��x��Jo���v�S���lI�&����rĚI�WH`��y���\̩w�K�3����~d��A� ����F��X1Q������4ڋ�霌�x,]i�|E=L7js�8v|ZN�@��&F�t?ʐ�V����j!������sh���O��lM ��U�G�*;/�To��ﭡ��=���������@;�<1�� ��ځhJ��P,\#�����G��C�����d�������;�|������~	͆�B^��̴fW]^�T��/٠�k�T?���8֮D���_cV]�pt;�JV��s�o����Fc2���Юh塑�ذqu\r�X9V������P\��;�ŉ�v�����q�<�疴6z�T�˱nݪظ����.p���
l��K�/jN[��u�S��8vtJ���To!sJ���/�P���5���r�c�ʕ1>:s3G��c��V�{ߣq��	�I�9����i<f�jT6{ ��W.��_=�R5v����L�}��J��+@�P���0s��"f
@Z~b��ӏƺ���������Ǟ�������-ٯ|�ݔƓF� k:�)�B���볝8��@4e��Z/1�?�3������h4�b瞣ی+��~y@�j�C����L�u~��Q˩eᡢ�ݐ�1فC�4�«� 1T����1ЭG�=���j�s�A�.s�>/�j�:�P�/(nnJ���(��P����S��G�k2��,���q�!��v��G33�U�t�ю�΂7��;K�ވڼL���X5��m['�c�l�cR��P���vP&Sd A��|��j�(�Kߡ���-�d^�у�o�s�-�����+7j������5��N�5�%�9QcG�]�NS�C3Jh,JMN�:q��IW�4X�U�B��į�j�/�J����:t���>�$}*jG&D�G�E=��E�P���s���oRM����n�h��`i��!i�ј\1��cdT�Ϧ��|��G��\M���C����h)֯���W�<n>+VǊ��j���g�o��zl�� ������|Sy.�3�17���ڦ{]ǌ�;��J}�j��8���إ Z2�%K�u|b,�ժ�\���N��챂d�Nv��^�.-}������, �B���ۑ��S��^[#�����Ğ�C�a�@������sq�бh��b\l|(�SS�Ly���(�ă���4
v�DS��Z#��Ż�рGfKx�%��C&J�9g�38:��VA`���HT�Q�D�L	V�1����x:��������\����E#�+bd|R��pK#��F�ތ~�kY=DU��N�4�G�Lec��a�G�&��ɼ����E���(J�6���ߍc{�����bs6f��2�ƆbL����P�%��4r.FTê��ʎ�_,20�}����c@&ΐ���=�;ܲ|�h�ı����[���1  T�<�`t^�fU��VcH����R��1��؈l<����ܜ4g�4*o�n�K�SU�s2O��NѤt���QD�1Bg�@�M
Bv�k�W�Զ�6��2;�?oJ/��g7M���B>׉��1.TF>�J��n�\e��Rf��Axp9Jʗi�����,�{=��dU�����V�84>��w��M���Ĵ��<n/W4��A�)	P#c�rŰ�2��x�!�Z1)�?��[���8M�1��c�jY���96>����˃����1�3�VQ>�b9�ؾ%~�߿�3G�[ O?�w���fǛ6���MwZ�u��.7�ݵ��?$�{vT�-�eS��2���-4Җ�:h+���$���uhD_�\F�@��A�L��=�Rr�MU�UU.�R3���b4d�.�(_�Ъā�5�*Mz�#ܪ!����c3�C�F�p̪˞S����\U&��+�V4�\������j4r�C�GD[VO��-t� O�A�ͷ��ə8x��lA�M����.�,R p���Jn��_H:mu+�q.��V���y���#|�����z�,u?�_�I�r[F�y�#&*��3�����kc�����,���?���oP����«�ƖuCq���]�m�Z]�z�n�b��Ҡ�k�,�LtU)بt�~1QZB�t?x"�2��K15׉��Ҭhwa���iAu�|�ՍWdN���GK\�6ろ+m�t��������� �o���gn��#�▻�K����dS9�����}��5�kt4�!-4d������M���{�y���q�7Nĳ.�˷�⟿�+v�S����`C��BlZ;/m^@���m��i�<m[��47.Y� 7�vۆјf1O1.��B��u������iCS�!!1��7Y��`W.K>�e�2�İ4�̞j�?�|ǎ�Me[�:i퇞8��-o������s�-�	q�H\�����ږ.����*��12�"6m9/�&�Iӭ���Pd+M������dTF&�:�.opT��[�*�FWǰ�׎(7��v��;[�qi�ёj�9t<蘑�1}���`-��?�>~$N>e��M2'�e��u���ػ{W;�7jSl��4��ND��ݱy�%QVy�8�wg�O������Xl��8P��W��=��=��7�:槎ǣ��S���X�q��7b���1�Z���=[��ꖭ[-���'����>&�{^�;����h4N�E^"��t����Q[���89�R��bC�ܻ�'R���S���P�vw@�O6�К[��S��<[��}��ص�`<�9ψ��-���=��ay#s�gXrH84�J6�X��G���[THyMHc�D�ƖT��=63�Nĉ��T�'�6ͣS�E�Ӧ���Q��0J��ctͶذeml�L��	�y*�)@�����Ǣ1�7f�����<��u��~�j��G�c�4�v�}_�]O���ػ�D�z��q���Wˡ�*L��i;�wz.������[o�}����VŬz��<�멘:vH��]6�U�;2��N�#s�)�G�m��.-����x� ��\*If�1�X���V:>;U�}��E�3kW�bͺ�X�au�^�>Vn�+6m�U>��ʕ����u��c���q|jV��׭���X�y�d�<��4�[ 'K �2c�)�����q��N<��S��5��(��M��r�5�i����l∑�\���ˌ��%����L
����ѹ�8Z�=ӕ�yX�H���Ҏ���m[��X�l[��y��1�S�ʒM>aЮM�Q����;�{o�{��qL�.{�z�1->	��.�&e�'��=;��g
q�=;�o�)��?��%o>0�/J������"�zr~!�iA�(c�D6�����Ÿ��cq�#�e���];����-ߌUk'br�EQ�(�<�e)�Ҹ�m��WEi`U���+�oV/UVa�2���ӱ�x.:<����ez��4>�ܲ�'�����u�m��2ɣGN�#=�{8�;��_f���dyc~*��d��X���(�G�:�ژF��Q���e<�P�w6T��\<���q˭���={�G���e4?��˟���^5矿=&�Fb`H2ٜ'�����+m���d@�v��CUvP�̢T�m���Ux��{�h��^�d1�g�)M)�2��?�P�!�1f
d�����ڵkdK��G�F=b{�o�h0�h*_5�OM�Ɓ�{��ǇeǪ��N�Y�2�VlP���� ܀����:��9,ᕪC��`�;�|�wG|��I�?3'Iv�x����O7!�Z�T�Ҕ�՞�p��?�3��1{PBE
���Ybr��@�nL�f?�� M�J� �
�������s
[�&S��h����7���4h�U���Ц���P�bРL�RL?J���-v���3�n[�E�c���S^f=��l R�I�Bf��_��;��`�g�������7�Ԙ���rE�R��p�8������`_7o�*U��<Ȩ�OG�H��{�W�hC�c����09��g��5X��4�[]![�ْ�����'w���Ѭ�ԭ���ܘ>�e0���%D�e&�cS���Y®�fT`[�Y�0�'�cY������Y9�U
5RX�'M��YU0�(т"������'n^ݰA��e��0$m�t�4�@lM�0k'x����+Ǥ 8)�+ǖ�b��5��X=	0���#k������S��B��br��2���1�qJ; �h���hC���?�+P.�_eYhEK��_���,*[�_f٩l�΢RԨ$[lzz~d(VH���N��	r�mf�l{�
���+{�~��, �`$0�z�O�4� �>B�x�CU�:�:ӿH-\x�<Ç��5��+Uԭk���%s�Ď�l�n�dS��`[��%TW���,�Y��x�>l``T��X5Z�.^W]�=�~�E��k.��^sq��y���%.�8$��D��bp�$�[�J���j��a,^x��x����������6�/[Wn�e&�*�FlakI��$s�mP�V�G�*[������U�*���2���v)�$�)HbUِo���w������,�$���E�!M�G��dL},�p$�s�-Ki�_�R	�"i�5H�FM��/DJȈ�RФh��C��x���ԐҲ��Kk��u%i*�A ����]hY%��!�n�U~%�*�ʋ��Q2#4��|�������~�`���Hܲo<�<2���ȍn�/�P�:K@����ʋ�C$a~�$��^��cO���W�,��"�\�_�"F������{��hx�mO�y���Aa�!#�j[[Rk�R���_#qҁ����d�2I���Zj�o[�0���%^���!�%κC;�
���^����箍�����A7��g���.r�J%��@�
��b��֡x�H6�s��^k&��a�H��R%P��<i�r)-d?
F�بt�h
�pu`0f�O�cw���q�-_�n�j<t�-qd����]Q]�<.�8k�!�P��]95݈��w�c߸'����ƭ����xg�z�]���c���1�P�ӎ��GV� ӯ�}tx@�KiZ���K&<ǸB�V����a4w{1j��8rl��=0��'��4�>*����R!j��8p�WJ��_v�dzѦ���+�Ŷ�#Q�e#�s�-��_#RmT�����*�����+_�¸���.�	�'NN1�R%�]I��U�F�{g N��1�@�P�_��P��^=�֯��������-�F=(���P��yj����*�x�P�X�/�+���-��;�cmi:*1��tfU�E���+Gb��D�Ԡo�h)V��a�U4��Tt�G�<�7J��ѭid��U;����;�_]�{!�ƅZ"�V��1��C6 ,*~��U4�+��U�N�ڷ7�Oգ�+G���d�������lQ��T��=G��31Y���p>֯���/�˯y�?��5V.�[ ��j�ti�J�͏Eԥ9f�ʫThit/ ���ǟ��ꑫI���.��8�N��e��Ǳ�G�A�nk~�z�1��ꑡX1���4��~�֒�<<:+G������������biX�n�+�֯*Ŀ}���%ϙ���}���j��ը��j�&b��ј\�ƳbB�Tٯ�s��B�����[K1*��w�Q�G��X�2 ��Y�Sq�z�_%R�e�
KE���2�.���ذ��S�[/�.�(֬�����؃Ń��G�;�u�����᝵����q���C;���ؾ9�.Z�ׯ��V�� �T���m� �"s���q��۶��]Ai���Ć��	H�V�[�w�A �D��/��:S������l�?��|7�������v�
��Scq�)����b�m�r��X�n�!� ���ϵV)��kblb� <h@x	�~ ��J���R�W\~Y̏�46>?Vm�*�E��Է�&m= ������ȄW��ɾ�@K��������~:6]|Yl�:��B`�#_���d�e?/�Qx��p�fOa��uK��A�j䗞�.��J��V�0�MP�18��uR�h6�����c�cwđ�w��]�Ǳ�o�C��'����]J�PO5�k�˼��}��[�<�&����y�}bL#�s�-�K����c�+�����������Kw����B����FEZ�.hH�����?�+��٣{b��ޘ9�;�:b~����U��F#�e��VD�<�������{\�>�J�H���������>�?�K�+����yB�Z"Z��5��x�H\yɖx���+7��vb~^ V�웛���7(���
p�A/P�����Z1<�"n��Gcc"���#�E���%� ӆ"*��rod"<�����8�������a[y|C��cN������;Չ��}qt�?�����-F]�W�b��'Z��U�W�0�Y�}袸"Z�!7��b%�5�'p��mĽ������ڴ������Inb�X�?v<�>�7v=��������b��m��5�,2g�4�c	Y T���2�����r�KCZ����6�(K+���x<��v����CGc��i��Ts�<Fƌ��`e1F����g<#�G��������|�OΎ9�n1���ƽ��{v>*>�TY��.�B ]�ht���5�@�W������ⲫ.��o�#��Xh�bbR�����k7Dm��B�yu�,����3����SqDÁ�����f0�x)����8z�d�7����\<��H<�؁xd��عc_�?p��Ç����q��L��q��t;6ǧk15ӎC'ڱ�`#����'��;���َ���[�_|��؝KnY�S.9i����/�������+NĦ�{�6�4�ty�A���S�)�bS ��.K�u�1{찧�FWnF[������<��Ӿ-/+�b�j �i���޸9���W�א�m.&W�a����٘���;�5���7������ص��Җ���S�G~<��Rwϓ.��4��,oF?���Q雍�����ӱ{ϡ���QU�_1/{�����y�8ȴ���l���=������@�D�]�,�2�4��8 s��e#���1M��O��l5$z�[>��ԙ����b�rX\��DO���X?�/~ɋ�E?�Q��9��=ǣ��I	;��;�f�ؕ�0��D���p�x�4U����Sq]sw�0yі��\?�>b��Ѩ�N�Q��Uq`߁8thVf6n��8�����yE\�����9�42(������ػ�� �Vב�w���zj���kS�^~E\w�1/��nB-#�#��W�$NH��\�Ƕ͛bX ��<�����	/�R�}��9��$��,R�zuȖ8h�|}*=�8���-��(���h�G�8�sѝ >G\�6+sc�5�؊�8����axf&n��c1^�����*���h5�T����{~H����� N3l��C����Bl�z~<r�m����F��#m����/��8v�.^i�aLc�����5�ը���'wn6�es�j�dB�E�k`�h�o6�����+��t[��Kd�_��-���y]=6'{��A�����PZ���q�Z~ &�{v����Xu�e�f����hh (j��6�v\z��Q�uO���]/JЂ�f�#Y^]��1������v���Xi�R����3,�b�6<3��.�Ҏk�"u�+�ncn�|Vl�;�Q�X��v^L�]��0�\h`���,7�ﺧv��i�/�p<ao�[�9�K��E�B� Lw�.���y<��*�Y{��g��S�D�o�2��!�/*�S{��<?�/6)+��:e���{z�]�4�V��˳67��=�w찶��f�W��|k�#��<��4����`'{ݱx�Х�\�P��"r�f�h��,5�?19.{Y����X�ai`�]�d�] �����3wP��4  � �V�V�����#jNik��럺6=����`f��,��Vt|�P���cx�&��uO�"�?��,��'A    IEND�B`�PK   U�tWJ1�~       jsons/user_defined.json��]o� ����ubq ;w�"M��jZ��)��A2$<l�����A�,�\�z������@+4���h�V*Ѡz��Z�8�	ؑ~������?n����l�;}��}ז�;jg�� v���l�߭͢_Л��]CxYU�fˢ����9�͒7yU�t�p�,��:/]f��E_�'��_d�O:���:�n�V�����etkw� O8a��.߾�'��	�8e'��\F%�ւ�i�#-����{�~���<�p��I�HR�� ������筶e%܂��kt\��� �f��l�H>	����_|F�x��H��y�̏�"�=�^|��H����,��"���y �b�g^|���L$p����#7@����r���p��<aS���E0��T �F��<eS��*�A0��D �N`��<jS��R��<�[- p�<O����<���ĥ�,�y��[x��A^y��"i/?|ͱe�o?X����}�����y��O��4�;<�!�;a�ܤ�F����v�9�PK
   U�tWm扴u  �                  cirkitFile.jsonPK
   �rmW�\>& %& /             �  images/27abb4c4-9cc3-40d1-807d-7d8b935f4094.pngPK
   U�tWJ1�~                 -> jsons/user_defined.jsonPK      �   w@   